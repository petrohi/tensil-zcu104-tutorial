module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_opcode,
  input  [3:0]  io_enq_bits_flags,
  input  [63:0] io_enq_bits_arguments,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_opcode,
  output [3:0]  io_deq_bits_flags,
  output [63:0] io_deq_bits_arguments
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_flags [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_flags_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_flags_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_flags_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_flags_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_flags_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_flags_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_flags_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_arguments [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_arguments_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_arguments_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_arguments_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_arguments_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_arguments_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_arguments_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_arguments_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_flags_io_deq_bits_MPORT_en = 1'h1;
  assign ram_flags_io_deq_bits_MPORT_addr = value_1;
  assign ram_flags_io_deq_bits_MPORT_data = ram_flags[ram_flags_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_flags_MPORT_data = io_enq_bits_flags;
  assign ram_flags_MPORT_addr = value;
  assign ram_flags_MPORT_mask = 1'h1;
  assign ram_flags_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_arguments_io_deq_bits_MPORT_en = 1'h1;
  assign ram_arguments_io_deq_bits_MPORT_addr = value_1;
  assign ram_arguments_io_deq_bits_MPORT_data = ram_arguments[ram_arguments_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_arguments_MPORT_data = io_enq_bits_arguments;
  assign ram_arguments_MPORT_addr = value;
  assign ram_arguments_MPORT_mask = 1'h1;
  assign ram_arguments_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_flags = ram_flags_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_arguments = ram_arguments_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_flags_MPORT_en & ram_flags_MPORT_mask) begin
      ram_flags[ram_flags_MPORT_addr] <= ram_flags_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_arguments_MPORT_en & ram_arguments_MPORT_mask) begin
      ram_arguments[ram_arguments_MPORT_addr] <= ram_arguments_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      value <= value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      value_1 <= value_1 + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_flags[initvar] = _RAND_1[3:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_arguments[initvar] = _RAND_2[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Counter(
  input         clock,
  input         reset,
  input         io_value_ready,
  output [20:0] io_value_bits,
  input         io_resetValue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] value; // @[Counter.scala 16:22]
  wire [20:0] _value_T_1 = value + 21'h1; // @[Counter.scala 24:22]
  assign io_value_bits = value; // @[Counter.scala 18:17]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 16:22]
      value <= 21'h0; // @[Counter.scala 16:22]
    end else if (io_resetValue) begin // @[Counter.scala 27:23]
      value <= 21'h0; // @[Counter.scala 28:11]
    end else if (io_value_ready) begin // @[Counter.scala 20:24]
      if (value == 21'h1fffff) begin // @[Counter.scala 21:31]
        value <= 21'h0; // @[Counter.scala 22:13]
      end else begin
        value <= _value_T_1; // @[Counter.scala 24:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[20:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CountBy(
  input         clock,
  input         reset,
  input         io_value_ready,
  output [20:0] io_value_bits,
  input  [20:0] io_step,
  input         io_resetValue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] value; // @[CountBy.scala 17:22]
  wire [21:0] _GEN_3 = {{1'd0}, io_step}; // @[CountBy.scala 22:24]
  wire [21:0] _T_1 = 22'h200000 - _GEN_3; // @[CountBy.scala 22:24]
  wire [21:0] _GEN_4 = {{1'd0}, value}; // @[CountBy.scala 22:16]
  wire [20:0] _value_T_1 = value + io_step; // @[CountBy.scala 25:22]
  assign io_value_bits = value; // @[CountBy.scala 19:17]
  always @(posedge clock) begin
    if (reset) begin // @[CountBy.scala 17:22]
      value <= 21'h0; // @[CountBy.scala 17:22]
    end else if (io_resetValue) begin // @[CountBy.scala 28:23]
      value <= 21'h0; // @[CountBy.scala 29:11]
    end else if (io_value_ready) begin // @[CountBy.scala 21:24]
      if (_GEN_4 >= _T_1) begin // @[CountBy.scala 22:36]
        value <= 21'h0; // @[CountBy.scala 23:13]
      end else begin
        value <= _value_T_1; // @[CountBy.scala 25:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[20:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SizeAndStrideHandler(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_write,
  input  [20:0] io_in_bits_address,
  input  [20:0] io_in_bits_size,
  input  [2:0]  io_in_bits_stride,
  input         io_in_bits_reverse,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_write,
  output [20:0] io_out_bits_address
);
  wire  sizeCounter_clock; // @[Counter.scala 34:19]
  wire  sizeCounter_reset; // @[Counter.scala 34:19]
  wire  sizeCounter_io_value_ready; // @[Counter.scala 34:19]
  wire [20:0] sizeCounter_io_value_bits; // @[Counter.scala 34:19]
  wire  sizeCounter_io_resetValue; // @[Counter.scala 34:19]
  wire  addressCounter_clock; // @[CountBy.scala 35:19]
  wire  addressCounter_reset; // @[CountBy.scala 35:19]
  wire  addressCounter_io_value_ready; // @[CountBy.scala 35:19]
  wire [20:0] addressCounter_io_value_bits; // @[CountBy.scala 35:19]
  wire [20:0] addressCounter_io_step; // @[CountBy.scala 35:19]
  wire  addressCounter_io_resetValue; // @[CountBy.scala 35:19]
  wire [7:0] stride = 8'h1 << io_in_bits_stride; // @[SizeAndStrideHandler.scala 30:20]
  wire [20:0] _io_out_bits_address_T_1 = io_in_bits_address - addressCounter_io_value_bits; // @[SizeAndStrideHandler.scala 46:44]
  wire [20:0] _io_out_bits_address_T_3 = io_in_bits_address + addressCounter_io_value_bits; // @[SizeAndStrideHandler.scala 48:44]
  wire  fire = io_in_valid & io_out_ready; // @[SizeAndStrideHandler.scala 51:23]
  Counter sizeCounter ( // @[Counter.scala 34:19]
    .clock(sizeCounter_clock),
    .reset(sizeCounter_reset),
    .io_value_ready(sizeCounter_io_value_ready),
    .io_value_bits(sizeCounter_io_value_bits),
    .io_resetValue(sizeCounter_io_resetValue)
  );
  CountBy addressCounter ( // @[CountBy.scala 35:19]
    .clock(addressCounter_clock),
    .reset(addressCounter_reset),
    .io_value_ready(addressCounter_io_value_ready),
    .io_value_bits(addressCounter_io_value_bits),
    .io_step(addressCounter_io_step),
    .io_resetValue(addressCounter_io_resetValue)
  );
  assign io_in_ready = sizeCounter_io_value_bits == io_in_bits_size & io_out_ready; // @[SizeAndStrideHandler.scala 53:52 54:14 58:14]
  assign io_out_valid = io_in_valid; // @[SizeAndStrideHandler.scala 35:16]
  assign io_out_bits_write = io_in_bits_write; // @[SizeAndStrideHandler.scala 38:34]
  assign io_out_bits_address = io_in_bits_reverse ? _io_out_bits_address_T_1 : _io_out_bits_address_T_3; // @[SizeAndStrideHandler.scala 45:25 46:25 48:25]
  assign sizeCounter_clock = clock;
  assign sizeCounter_reset = reset;
  assign sizeCounter_io_value_ready = sizeCounter_io_value_bits == io_in_bits_size ? 1'h0 : fire; // @[Counter.scala 36:22 SizeAndStrideHandler.scala 53:52 59:32]
  assign sizeCounter_io_resetValue = sizeCounter_io_value_bits == io_in_bits_size & fire; // @[Counter.scala 35:21 SizeAndStrideHandler.scala 53:52 55:31]
  assign addressCounter_clock = clock;
  assign addressCounter_reset = reset;
  assign addressCounter_io_value_ready = sizeCounter_io_value_bits == io_in_bits_size ? 1'h0 : fire; // @[Counter.scala 36:22 SizeAndStrideHandler.scala 53:52 59:32]
  assign addressCounter_io_step = {{13'd0}, stride}; // @[CountBy.scala 36:15]
  assign addressCounter_io_resetValue = sizeCounter_io_value_bits == io_in_bits_size & fire; // @[Counter.scala 35:21 SizeAndStrideHandler.scala 53:52 55:31]
endmodule
module StrideHandler(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_write,
  input  [20:0] io_in_bits_address,
  input  [20:0] io_in_bits_size,
  input  [2:0]  io_in_bits_stride,
  input         io_in_bits_reverse,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_write,
  output [20:0] io_out_bits_address,
  output [20:0] io_out_bits_size
);
  wire  handler_clock; // @[StrideHandler.scala 27:23]
  wire  handler_reset; // @[StrideHandler.scala 27:23]
  wire  handler_io_in_ready; // @[StrideHandler.scala 27:23]
  wire  handler_io_in_valid; // @[StrideHandler.scala 27:23]
  wire  handler_io_in_bits_write; // @[StrideHandler.scala 27:23]
  wire [20:0] handler_io_in_bits_address; // @[StrideHandler.scala 27:23]
  wire [20:0] handler_io_in_bits_size; // @[StrideHandler.scala 27:23]
  wire [2:0] handler_io_in_bits_stride; // @[StrideHandler.scala 27:23]
  wire  handler_io_in_bits_reverse; // @[StrideHandler.scala 27:23]
  wire  handler_io_out_ready; // @[StrideHandler.scala 27:23]
  wire  handler_io_out_valid; // @[StrideHandler.scala 27:23]
  wire  handler_io_out_bits_write; // @[StrideHandler.scala 27:23]
  wire [20:0] handler_io_out_bits_address; // @[StrideHandler.scala 27:23]
  SizeAndStrideHandler handler ( // @[StrideHandler.scala 27:23]
    .clock(handler_clock),
    .reset(handler_reset),
    .io_in_ready(handler_io_in_ready),
    .io_in_valid(handler_io_in_valid),
    .io_in_bits_write(handler_io_in_bits_write),
    .io_in_bits_address(handler_io_in_bits_address),
    .io_in_bits_size(handler_io_in_bits_size),
    .io_in_bits_stride(handler_io_in_bits_stride),
    .io_in_bits_reverse(handler_io_in_bits_reverse),
    .io_out_ready(handler_io_out_ready),
    .io_out_valid(handler_io_out_valid),
    .io_out_bits_write(handler_io_out_bits_write),
    .io_out_bits_address(handler_io_out_bits_address)
  );
  assign io_in_ready = io_in_bits_stride == 3'h0 ? io_out_ready : handler_io_in_ready; // @[StrideHandler.scala 41:32 49:14 52:19]
  assign io_out_valid = io_in_bits_stride == 3'h0 ? io_in_valid : handler_io_out_valid; // @[StrideHandler.scala 41:32 50:18 61:18]
  assign io_out_bits_write = io_in_bits_stride == 3'h0 ? io_in_bits_write : handler_io_out_bits_write; // @[StrideHandler.scala 41:32 44:36 55:36]
  assign io_out_bits_address = io_in_bits_stride == 3'h0 ? io_in_bits_address : handler_io_out_bits_address; // @[StrideHandler.scala 41:32 47:25 58:25]
  assign io_out_bits_size = io_in_bits_stride == 3'h0 ? io_in_bits_size : 21'h0; // @[StrideHandler.scala 41:32 48:22 59:22]
  assign handler_clock = clock;
  assign handler_reset = reset;
  assign handler_io_in_valid = io_in_bits_stride == 3'h0 ? 1'h0 : io_in_valid; // @[StrideHandler.scala 37:23 41:32 52:19]
  assign handler_io_in_bits_write = io_in_bits_stride == 3'h0 ? 1'h0 : io_in_bits_write; // @[StrideHandler.scala 38:22 41:32 52:19]
  assign handler_io_in_bits_address = io_in_bits_stride == 3'h0 ? 21'h0 : io_in_bits_address; // @[StrideHandler.scala 38:22 41:32 52:19]
  assign handler_io_in_bits_size = io_in_bits_stride == 3'h0 ? 21'h0 : io_in_bits_size; // @[StrideHandler.scala 38:22 41:32 52:19]
  assign handler_io_in_bits_stride = io_in_bits_stride == 3'h0 ? 3'h0 : io_in_bits_stride; // @[StrideHandler.scala 38:22 41:32 52:19]
  assign handler_io_in_bits_reverse = io_in_bits_stride == 3'h0 ? 1'h0 : io_in_bits_reverse; // @[StrideHandler.scala 38:22 41:32 52:19]
  assign handler_io_out_ready = io_in_bits_stride == 3'h0 ? 1'h0 : io_out_ready; // @[StrideHandler.scala 39:24 41:32 60:26]
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_write,
  input  [20:0] io_enq_bits_address,
  input  [20:0] io_enq_bits_size,
  input  [2:0]  io_enq_bits_stride,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_write,
  output [20:0] io_deq_bits_address,
  output [20:0] io_deq_bits_size,
  output [2:0]  io_deq_bits_stride,
  output        io_deq_bits_reverse
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  ram_write [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_en; // @[Decoupled.scala 259:95]
  reg [20:0] ram_address [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [20:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [20:0] ram_address_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 259:95]
  reg [20:0] ram_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [20:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [20:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_stride [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_stride_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_stride_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_stride_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_stride_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_stride_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_stride_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_stride_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_reverse [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_reverse_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_reverse_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_reverse_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_reverse_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_reverse_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_reverse_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_reverse_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_13 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_13 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_write_io_deq_bits_MPORT_en = 1'h1;
  assign ram_write_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_write_io_deq_bits_MPORT_data = ram_write[ram_write_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_write_MPORT_data = io_enq_bits_write;
  assign ram_write_MPORT_addr = 1'h0;
  assign ram_write_MPORT_mask = 1'h1;
  assign ram_write_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = 1'h0;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign ram_stride_io_deq_bits_MPORT_en = 1'h1;
  assign ram_stride_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_stride_io_deq_bits_MPORT_data = ram_stride[ram_stride_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_stride_MPORT_data = io_enq_bits_stride;
  assign ram_stride_MPORT_addr = 1'h0;
  assign ram_stride_MPORT_mask = 1'h1;
  assign ram_stride_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign ram_reverse_io_deq_bits_MPORT_en = 1'h1;
  assign ram_reverse_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_reverse_io_deq_bits_MPORT_data = ram_reverse[ram_reverse_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_reverse_MPORT_data = 1'h0;
  assign ram_reverse_MPORT_addr = 1'h0;
  assign ram_reverse_MPORT_mask = 1'h1;
  assign ram_reverse_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_write = empty ? io_enq_bits_write : ram_write_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_address = empty ? io_enq_bits_address : ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_stride = empty ? io_enq_bits_stride : ram_stride_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_reverse = empty ? 1'h0 : ram_reverse_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_write_MPORT_en & ram_write_MPORT_mask) begin
      ram_write[ram_write_MPORT_addr] <= ram_write_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_stride_MPORT_en & ram_stride_MPORT_mask) begin
      ram_stride[ram_stride_MPORT_addr] <= ram_stride_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_reverse_MPORT_en & ram_reverse_MPORT_mask) begin
      ram_reverse[ram_reverse_MPORT_addr] <= ram_reverse_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_write[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_address[initvar] = _RAND_1[20:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[20:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_stride[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_reverse[initvar] = _RAND_4[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Counter_2(
  input         clock,
  input         reset,
  input         io_value_ready,
  output [13:0] io_value_bits,
  input         io_resetValue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [13:0] value; // @[Counter.scala 16:22]
  wire [13:0] _value_T_1 = value + 14'h1; // @[Counter.scala 24:22]
  assign io_value_bits = value; // @[Counter.scala 18:17]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 16:22]
      value <= 14'h0; // @[Counter.scala 16:22]
    end else if (io_resetValue) begin // @[Counter.scala 27:23]
      value <= 14'h0; // @[Counter.scala 28:11]
    end else if (io_value_ready) begin // @[Counter.scala 20:24]
      if (value == 14'h3fff) begin // @[Counter.scala 21:31]
        value <= 14'h0; // @[Counter.scala 22:13]
      end else begin
        value <= _value_T_1; // @[Counter.scala 24:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[13:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CountBy_2(
  input         clock,
  input         reset,
  input         io_value_ready,
  output [13:0] io_value_bits,
  input  [13:0] io_step,
  input         io_resetValue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [13:0] value; // @[CountBy.scala 17:22]
  wire [14:0] _GEN_3 = {{1'd0}, io_step}; // @[CountBy.scala 22:24]
  wire [14:0] _T_1 = 15'h4000 - _GEN_3; // @[CountBy.scala 22:24]
  wire [14:0] _GEN_4 = {{1'd0}, value}; // @[CountBy.scala 22:16]
  wire [13:0] _value_T_1 = value + io_step; // @[CountBy.scala 25:22]
  assign io_value_bits = value; // @[CountBy.scala 19:17]
  always @(posedge clock) begin
    if (reset) begin // @[CountBy.scala 17:22]
      value <= 14'h0; // @[CountBy.scala 17:22]
    end else if (io_resetValue) begin // @[CountBy.scala 28:23]
      value <= 14'h0; // @[CountBy.scala 29:11]
    end else if (io_value_ready) begin // @[CountBy.scala 21:24]
      if (_GEN_4 >= _T_1) begin // @[CountBy.scala 22:36]
        value <= 14'h0; // @[CountBy.scala 23:13]
      end else begin
        value <= _value_T_1; // @[CountBy.scala 25:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[13:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SizeAndStrideHandler_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_write,
  input  [13:0] io_in_bits_address,
  input  [13:0] io_in_bits_size,
  input  [2:0]  io_in_bits_stride,
  input         io_in_bits_reverse,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_write,
  output [13:0] io_out_bits_address
);
  wire  sizeCounter_clock; // @[Counter.scala 34:19]
  wire  sizeCounter_reset; // @[Counter.scala 34:19]
  wire  sizeCounter_io_value_ready; // @[Counter.scala 34:19]
  wire [13:0] sizeCounter_io_value_bits; // @[Counter.scala 34:19]
  wire  sizeCounter_io_resetValue; // @[Counter.scala 34:19]
  wire  addressCounter_clock; // @[CountBy.scala 35:19]
  wire  addressCounter_reset; // @[CountBy.scala 35:19]
  wire  addressCounter_io_value_ready; // @[CountBy.scala 35:19]
  wire [13:0] addressCounter_io_value_bits; // @[CountBy.scala 35:19]
  wire [13:0] addressCounter_io_step; // @[CountBy.scala 35:19]
  wire  addressCounter_io_resetValue; // @[CountBy.scala 35:19]
  wire [7:0] stride = 8'h1 << io_in_bits_stride; // @[SizeAndStrideHandler.scala 30:20]
  wire [13:0] _io_out_bits_address_T_1 = io_in_bits_address - addressCounter_io_value_bits; // @[SizeAndStrideHandler.scala 46:44]
  wire [13:0] _io_out_bits_address_T_3 = io_in_bits_address + addressCounter_io_value_bits; // @[SizeAndStrideHandler.scala 48:44]
  wire  fire = io_in_valid & io_out_ready; // @[SizeAndStrideHandler.scala 51:23]
  Counter_2 sizeCounter ( // @[Counter.scala 34:19]
    .clock(sizeCounter_clock),
    .reset(sizeCounter_reset),
    .io_value_ready(sizeCounter_io_value_ready),
    .io_value_bits(sizeCounter_io_value_bits),
    .io_resetValue(sizeCounter_io_resetValue)
  );
  CountBy_2 addressCounter ( // @[CountBy.scala 35:19]
    .clock(addressCounter_clock),
    .reset(addressCounter_reset),
    .io_value_ready(addressCounter_io_value_ready),
    .io_value_bits(addressCounter_io_value_bits),
    .io_step(addressCounter_io_step),
    .io_resetValue(addressCounter_io_resetValue)
  );
  assign io_in_ready = sizeCounter_io_value_bits == io_in_bits_size & io_out_ready; // @[SizeAndStrideHandler.scala 53:52 54:14 58:14]
  assign io_out_valid = io_in_valid; // @[SizeAndStrideHandler.scala 35:16]
  assign io_out_bits_write = io_in_bits_write; // @[SizeAndStrideHandler.scala 38:34]
  assign io_out_bits_address = io_in_bits_reverse ? _io_out_bits_address_T_1 : _io_out_bits_address_T_3; // @[SizeAndStrideHandler.scala 45:25 46:25 48:25]
  assign sizeCounter_clock = clock;
  assign sizeCounter_reset = reset;
  assign sizeCounter_io_value_ready = sizeCounter_io_value_bits == io_in_bits_size ? 1'h0 : fire; // @[Counter.scala 36:22 SizeAndStrideHandler.scala 53:52 59:32]
  assign sizeCounter_io_resetValue = sizeCounter_io_value_bits == io_in_bits_size & fire; // @[Counter.scala 35:21 SizeAndStrideHandler.scala 53:52 55:31]
  assign addressCounter_clock = clock;
  assign addressCounter_reset = reset;
  assign addressCounter_io_value_ready = sizeCounter_io_value_bits == io_in_bits_size ? 1'h0 : fire; // @[Counter.scala 36:22 SizeAndStrideHandler.scala 53:52 59:32]
  assign addressCounter_io_step = {{6'd0}, stride}; // @[CountBy.scala 36:15]
  assign addressCounter_io_resetValue = sizeCounter_io_value_bits == io_in_bits_size & fire; // @[Counter.scala 35:21 SizeAndStrideHandler.scala 53:52 55:31]
endmodule
module LockPool(
  input         clock,
  input         reset,
  output        io_actor_0_in_ready,
  input         io_actor_0_in_valid,
  input         io_actor_0_in_bits_write,
  input  [13:0] io_actor_0_in_bits_address,
  input  [13:0] io_actor_0_in_bits_size,
  input  [2:0]  io_actor_0_in_bits_stride,
  input         io_actor_0_in_bits_reverse,
  input         io_actor_0_out_ready,
  output        io_actor_0_out_valid,
  output        io_actor_0_out_bits_write,
  output [13:0] io_actor_0_out_bits_address,
  output [13:0] io_actor_0_out_bits_size,
  output [2:0]  io_actor_0_out_bits_stride,
  output        io_actor_0_out_bits_reverse,
  output        io_actor_1_in_ready,
  input         io_actor_1_in_valid,
  input         io_actor_1_in_bits_write,
  input  [13:0] io_actor_1_in_bits_address,
  input  [13:0] io_actor_1_in_bits_size,
  input  [2:0]  io_actor_1_in_bits_stride,
  input         io_actor_1_out_ready,
  output        io_actor_1_out_valid,
  output        io_actor_1_out_bits_write,
  output [13:0] io_actor_1_out_bits_address,
  output [13:0] io_actor_1_out_bits_size,
  output [2:0]  io_actor_1_out_bits_stride,
  output        io_actor_1_out_bits_reverse,
  output        io_lock_ready,
  input         io_lock_valid,
  input         io_lock_bits_cond_write,
  input  [13:0] io_lock_bits_cond_address,
  input  [13:0] io_lock_bits_cond_size,
  input  [2:0]  io_lock_bits_cond_stride,
  input         io_lock_bits_cond_reverse,
  input         io_lock_bits_lock,
  input         io_lock_bits_by
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg  lock_0_cond_write; // @[LockPool.scala 55:21]
  reg [13:0] lock_0_cond_address; // @[LockPool.scala 55:21]
  reg [13:0] lock_0_cond_size; // @[LockPool.scala 55:21]
  reg [2:0] lock_0_cond_stride; // @[LockPool.scala 55:21]
  reg  lock_0_cond_reverse; // @[LockPool.scala 55:21]
  reg  lock_0_held; // @[LockPool.scala 55:21]
  reg  lock_0_by; // @[LockPool.scala 55:21]
  reg  lock_1_cond_write; // @[LockPool.scala 55:21]
  reg [13:0] lock_1_cond_address; // @[LockPool.scala 55:21]
  reg [13:0] lock_1_cond_size; // @[LockPool.scala 55:21]
  reg [2:0] lock_1_cond_stride; // @[LockPool.scala 55:21]
  reg  lock_1_cond_reverse; // @[LockPool.scala 55:21]
  reg  lock_1_held; // @[LockPool.scala 55:21]
  reg  lock_1_by; // @[LockPool.scala 55:21]
  wire [13:0] block_requiredLockId = io_actor_0_in_bits_address / 14'h2000; // @[Decoder.scala 191:15]
  wire  _GEN_1 = block_requiredLockId[0] ? lock_1_by : lock_0_by; // @[LockPool.scala 70:{45,45}]
  wire  _GEN_3 = block_requiredLockId[0] ? lock_1_held : lock_0_held; // @[LockPool.scala 70:{26,26}]
  wire  _block_blocked_T_2 = io_lock_ready & io_lock_valid; // @[Decoupled.scala 50:35]
  wire [13:0] _GEN_224 = {{13'd0}, io_lock_bits_lock}; // @[LockPool.scala 70:101]
  wire  block_blocked = _GEN_3 & _GEN_1 | _block_blocked_T_2 & _GEN_224 == block_requiredLockId & io_lock_bits_by; // @[LockPool.scala 70:55]
  wire  _GEN_4 = ~block_blocked & io_actor_0_out_ready; // @[LockPool.scala 66:13 71:20 73:24]
  wire  _GEN_5 = ~block_blocked & io_actor_0_in_valid; // @[LockPool.scala 71:20 Decoupled.scala 72:20 LockPool.scala 73:24]
  wire [13:0] block_requiredLockId_1 = io_actor_1_in_bits_address / 14'h2000; // @[Decoder.scala 191:15]
  wire  _GEN_12 = block_requiredLockId_1[0] ? lock_1_by : lock_0_by; // @[LockPool.scala 70:{45,45}]
  wire  _GEN_14 = block_requiredLockId_1[0] ? lock_1_held : lock_0_held; // @[LockPool.scala 70:{26,26}]
  wire  block_blocked_1 = _GEN_14 & ~_GEN_12 | _block_blocked_T_2 & _GEN_224 == block_requiredLockId_1 & ~
    io_lock_bits_by; // @[LockPool.scala 70:55]
  wire  _GEN_15 = ~block_blocked_1 & io_actor_1_out_ready; // @[LockPool.scala 66:13 71:20 73:24]
  wire  _GEN_16 = ~block_blocked_1 & io_actor_1_in_valid; // @[LockPool.scala 71:20 Decoupled.scala 72:20 LockPool.scala 73:24]
  wire  _GEN_197 = lock_0_by ? io_actor_1_out_ready : io_actor_0_out_ready; // @[LockPool.scala 140:{32,32}]
  wire  _GEN_194 = ~lock_0_by ? _GEN_197 : _GEN_4; // @[LockPool.scala 140:{32,32}]
  wire  actor_0_ready = block_blocked & block_blocked_1 ? _GEN_194 : _GEN_4; // @[LockPool.scala 139:40]
  wire  _GEN_195 = lock_0_by ? _GEN_197 : _GEN_15; // @[LockPool.scala 140:{32,32}]
  wire  actor_1_ready = block_blocked & block_blocked_1 ? _GEN_195 : _GEN_15; // @[LockPool.scala 139:40]
  wire  _GEN_23 = io_lock_bits_by ? actor_1_ready : actor_0_ready; // @[Decoupled.scala 50:{35,35}]
  wire  _GEN_25 = io_lock_bits_by ? io_actor_1_in_valid : io_actor_0_in_valid; // @[Decoupled.scala 50:{35,35}]
  wire  _incomingObserved_T = _GEN_23 & _GEN_25; // @[Decoupled.scala 50:35]
  wire [13:0] _GEN_27 = io_lock_bits_by ? io_actor_1_in_bits_address : io_actor_0_in_bits_address; // @[MemControl.scala 21:{13,13}]
  wire  _GEN_29 = io_lock_bits_by ? io_actor_1_in_bits_write : io_actor_0_in_bits_write; // @[MemControl.scala 21:{40,40}]
  wire [13:0] _GEN_31 = io_lock_bits_by ? io_actor_1_in_bits_size : io_actor_0_in_bits_size; // @[MemControl.scala 21:{64,64}]
  wire [2:0] _GEN_33 = io_lock_bits_by ? io_actor_1_in_bits_stride : io_actor_0_in_bits_stride; // @[MemControl.scala 21:{89,89}]
  wire  _GEN_35 = io_lock_bits_by ? 1'h0 : io_actor_0_in_bits_reverse; // @[MemControl.scala 21:{117,117}]
  wire  _incomingObserved_T_10 = _GEN_27 == io_lock_bits_cond_address & _GEN_29 == io_lock_bits_cond_write & _GEN_31 ==
    io_lock_bits_cond_size & _GEN_33 == io_lock_bits_cond_stride & _GEN_35 == io_lock_bits_cond_reverse; // @[MemControl.scala 21:106]
  wire  incomingObserved = io_lock_valid & _incomingObserved_T & _incomingObserved_T_10; // @[LockPool.scala 98:58]
  wire  _GEN_37 = io_lock_bits_lock ? lock_1_by : lock_0_by; // @[LockPool.scala 104:{68,68}]
  wire  _GEN_39 = io_lock_bits_lock ? lock_1_held : lock_0_held; // @[LockPool.scala 104:{45,45}]
  wire  incoming = ~io_lock_bits_lock; // @[LockPool.scala 106:42]
  wire  _GEN_41 = lock_0_by ? actor_1_ready : actor_0_ready; // @[Decoupled.scala 50:{35,35}]
  wire  _GEN_43 = lock_0_by ? io_actor_1_in_valid : io_actor_0_in_valid; // @[Decoupled.scala 50:{35,35}]
  wire  _observed_T = _GEN_41 & _GEN_43; // @[Decoupled.scala 50:35]
  wire [13:0] _GEN_45 = lock_0_by ? io_actor_1_in_bits_address : io_actor_0_in_bits_address; // @[MemControl.scala 21:{13,13}]
  wire  _GEN_47 = lock_0_by ? io_actor_1_in_bits_write : io_actor_0_in_bits_write; // @[MemControl.scala 21:{40,40}]
  wire [13:0] _GEN_49 = lock_0_by ? io_actor_1_in_bits_size : io_actor_0_in_bits_size; // @[MemControl.scala 21:{64,64}]
  wire [2:0] _GEN_51 = lock_0_by ? io_actor_1_in_bits_stride : io_actor_0_in_bits_stride; // @[MemControl.scala 21:{89,89}]
  wire  _GEN_53 = lock_0_by ? 1'h0 : io_actor_0_in_bits_reverse; // @[MemControl.scala 21:{117,117}]
  wire  _observed_T_9 = _GEN_45 == lock_0_cond_address & _GEN_47 == lock_0_cond_write & _GEN_49 == lock_0_cond_size &
    _GEN_51 == lock_0_cond_stride & _GEN_53 == lock_0_cond_reverse; // @[MemControl.scala 21:106]
  wire  observed = _observed_T & _observed_T_9; // @[LockPool.scala 107:37]
  wire  _GEN_55 = io_lock_valid ? io_lock_bits_by : lock_0_by; // @[LockPool.scala 86:29 88:12 55:21]
  wire  _GEN_56 = io_lock_valid ? io_lock_bits_cond_write : lock_0_cond_write; // @[LockPool.scala 86:29 89:14 55:21]
  wire [13:0] _GEN_57 = io_lock_valid ? io_lock_bits_cond_address : lock_0_cond_address; // @[LockPool.scala 86:29 89:14 55:21]
  wire [13:0] _GEN_58 = io_lock_valid ? io_lock_bits_cond_size : lock_0_cond_size; // @[LockPool.scala 86:29 89:14 55:21]
  wire [2:0] _GEN_59 = io_lock_valid ? io_lock_bits_cond_stride : lock_0_cond_stride; // @[LockPool.scala 86:29 89:14 55:21]
  wire  _GEN_60 = io_lock_valid ? io_lock_bits_cond_reverse : lock_0_cond_reverse; // @[LockPool.scala 86:29 89:14 55:21]
  wire  _GEN_61 = incomingObserved ? 1'h0 : io_lock_valid; // @[LockPool.scala 111:34 93:12]
  wire  _GEN_62 = incomingObserved ? lock_0_by : _GEN_55; // @[LockPool.scala 111:34 55:21]
  wire  _GEN_63 = incomingObserved ? lock_0_cond_write : _GEN_56; // @[LockPool.scala 111:34 55:21]
  wire [13:0] _GEN_64 = incomingObserved ? lock_0_cond_address : _GEN_57; // @[LockPool.scala 111:34 55:21]
  wire [13:0] _GEN_65 = incomingObserved ? lock_0_cond_size : _GEN_58; // @[LockPool.scala 111:34 55:21]
  wire [2:0] _GEN_66 = incomingObserved ? lock_0_cond_stride : _GEN_59; // @[LockPool.scala 111:34 55:21]
  wire  _GEN_67 = incomingObserved ? lock_0_cond_reverse : _GEN_60; // @[LockPool.scala 111:34 55:21]
  wire  _GEN_68 = incoming & _GEN_61; // @[LockPool.scala 110:24 93:12]
  wire  _GEN_75 = io_lock_valid | lock_0_held; // @[LockPool.scala 86:29 87:14 55:21]
  wire  _GEN_76 = lock_0_by == io_lock_bits_by ? _GEN_75 : lock_0_held; // @[LockPool.scala 123:46 55:21]
  wire  _GEN_77 = lock_0_by == io_lock_bits_by ? _GEN_55 : lock_0_by; // @[LockPool.scala 123:46 55:21]
  wire  _GEN_78 = lock_0_by == io_lock_bits_by ? _GEN_56 : lock_0_cond_write; // @[LockPool.scala 123:46 55:21]
  wire [13:0] _GEN_79 = lock_0_by == io_lock_bits_by ? _GEN_57 : lock_0_cond_address; // @[LockPool.scala 123:46 55:21]
  wire [13:0] _GEN_80 = lock_0_by == io_lock_bits_by ? _GEN_58 : lock_0_cond_size; // @[LockPool.scala 123:46 55:21]
  wire [2:0] _GEN_81 = lock_0_by == io_lock_bits_by ? _GEN_59 : lock_0_cond_stride; // @[LockPool.scala 123:46 55:21]
  wire  _GEN_82 = lock_0_by == io_lock_bits_by ? _GEN_60 : lock_0_cond_reverse; // @[LockPool.scala 123:46 55:21]
  wire  _GEN_119 = lock_1_by ? actor_1_ready : actor_0_ready; // @[Decoupled.scala 50:{35,35}]
  wire  _GEN_121 = lock_1_by ? io_actor_1_in_valid : io_actor_0_in_valid; // @[Decoupled.scala 50:{35,35}]
  wire  _observed_T_10 = _GEN_119 & _GEN_121; // @[Decoupled.scala 50:35]
  wire [13:0] _GEN_123 = lock_1_by ? io_actor_1_in_bits_address : io_actor_0_in_bits_address; // @[MemControl.scala 21:{13,13}]
  wire  _GEN_125 = lock_1_by ? io_actor_1_in_bits_write : io_actor_0_in_bits_write; // @[MemControl.scala 21:{40,40}]
  wire [13:0] _GEN_127 = lock_1_by ? io_actor_1_in_bits_size : io_actor_0_in_bits_size; // @[MemControl.scala 21:{64,64}]
  wire [2:0] _GEN_129 = lock_1_by ? io_actor_1_in_bits_stride : io_actor_0_in_bits_stride; // @[MemControl.scala 21:{89,89}]
  wire  _GEN_131 = lock_1_by ? 1'h0 : io_actor_0_in_bits_reverse; // @[MemControl.scala 21:{117,117}]
  wire  _observed_T_19 = _GEN_123 == lock_1_cond_address & _GEN_125 == lock_1_cond_write & _GEN_127 == lock_1_cond_size
     & _GEN_129 == lock_1_cond_stride & _GEN_131 == lock_1_cond_reverse; // @[MemControl.scala 21:106]
  wire  observed_1 = _observed_T_10 & _observed_T_19; // @[LockPool.scala 107:37]
  wire  _GEN_132 = io_lock_valid ? io_lock_bits_by : lock_1_by; // @[LockPool.scala 86:29 88:12 55:21]
  wire  _GEN_133 = io_lock_valid ? io_lock_bits_cond_write : lock_1_cond_write; // @[LockPool.scala 86:29 89:14 55:21]
  wire [13:0] _GEN_134 = io_lock_valid ? io_lock_bits_cond_address : lock_1_cond_address; // @[LockPool.scala 86:29 89:14 55:21]
  wire [13:0] _GEN_135 = io_lock_valid ? io_lock_bits_cond_size : lock_1_cond_size; // @[LockPool.scala 86:29 89:14 55:21]
  wire [2:0] _GEN_136 = io_lock_valid ? io_lock_bits_cond_stride : lock_1_cond_stride; // @[LockPool.scala 86:29 89:14 55:21]
  wire  _GEN_137 = io_lock_valid ? io_lock_bits_cond_reverse : lock_1_cond_reverse; // @[LockPool.scala 86:29 89:14 55:21]
  wire  _GEN_138 = incomingObserved ? lock_1_by : _GEN_132; // @[LockPool.scala 111:34 55:21]
  wire  _GEN_139 = incomingObserved ? lock_1_cond_write : _GEN_133; // @[LockPool.scala 111:34 55:21]
  wire [13:0] _GEN_140 = incomingObserved ? lock_1_cond_address : _GEN_134; // @[LockPool.scala 111:34 55:21]
  wire [13:0] _GEN_141 = incomingObserved ? lock_1_cond_size : _GEN_135; // @[LockPool.scala 111:34 55:21]
  wire [2:0] _GEN_142 = incomingObserved ? lock_1_cond_stride : _GEN_136; // @[LockPool.scala 111:34 55:21]
  wire  _GEN_143 = incomingObserved ? lock_1_cond_reverse : _GEN_137; // @[LockPool.scala 111:34 55:21]
  wire  _GEN_144 = io_lock_bits_lock & _GEN_61; // @[LockPool.scala 110:24 93:12]
  wire  _GEN_151 = io_lock_valid | lock_1_held; // @[LockPool.scala 86:29 87:14 55:21]
  wire  _GEN_152 = lock_1_by == io_lock_bits_by ? _GEN_151 : lock_1_held; // @[LockPool.scala 123:46 55:21]
  wire  _GEN_153 = lock_1_by == io_lock_bits_by ? _GEN_132 : lock_1_by; // @[LockPool.scala 123:46 55:21]
  wire  _GEN_154 = lock_1_by == io_lock_bits_by ? _GEN_133 : lock_1_cond_write; // @[LockPool.scala 123:46 55:21]
  wire [13:0] _GEN_155 = lock_1_by == io_lock_bits_by ? _GEN_134 : lock_1_cond_address; // @[LockPool.scala 123:46 55:21]
  wire [13:0] _GEN_156 = lock_1_by == io_lock_bits_by ? _GEN_135 : lock_1_cond_size; // @[LockPool.scala 123:46 55:21]
  wire [2:0] _GEN_157 = lock_1_by == io_lock_bits_by ? _GEN_136 : lock_1_cond_stride; // @[LockPool.scala 123:46 55:21]
  wire  _GEN_158 = lock_1_by == io_lock_bits_by ? _GEN_137 : lock_1_cond_reverse; // @[LockPool.scala 123:46 55:21]
  wire  _GEN_198 = ~lock_0_by ? _GEN_43 : _GEN_5; // @[LockPool.scala 140:{32,32}]
  wire  _GEN_199 = lock_0_by ? _GEN_43 : _GEN_16; // @[LockPool.scala 140:{32,32}]
  wire  _GEN_200 = ~lock_0_by ? _GEN_47 : io_actor_0_in_bits_write; // @[LockPool.scala 140:{32,32}]
  wire  _GEN_201 = lock_0_by ? _GEN_47 : io_actor_1_in_bits_write; // @[LockPool.scala 140:{32,32}]
  wire [13:0] _GEN_202 = ~lock_0_by ? _GEN_45 : io_actor_0_in_bits_address; // @[LockPool.scala 140:{32,32}]
  wire [13:0] _GEN_203 = lock_0_by ? _GEN_45 : io_actor_1_in_bits_address; // @[LockPool.scala 140:{32,32}]
  wire [13:0] _GEN_204 = ~lock_0_by ? _GEN_49 : io_actor_0_in_bits_size; // @[LockPool.scala 140:{32,32}]
  wire [13:0] _GEN_205 = lock_0_by ? _GEN_49 : io_actor_1_in_bits_size; // @[LockPool.scala 140:{32,32}]
  wire [2:0] _GEN_206 = ~lock_0_by ? _GEN_51 : io_actor_0_in_bits_stride; // @[LockPool.scala 140:{32,32}]
  wire [2:0] _GEN_207 = lock_0_by ? _GEN_51 : io_actor_1_in_bits_stride; // @[LockPool.scala 140:{32,32}]
  wire  _GEN_208 = ~lock_0_by ? _GEN_53 : io_actor_0_in_bits_reverse; // @[LockPool.scala 140:{32,32}]
  wire  _GEN_209 = lock_0_by & _GEN_53; // @[LockPool.scala 140:{32,32}]
  assign io_actor_0_in_ready = block_blocked & block_blocked_1 ? _GEN_194 : _GEN_4; // @[LockPool.scala 139:40]
  assign io_actor_0_out_valid = block_blocked & block_blocked_1 ? _GEN_198 : _GEN_5; // @[LockPool.scala 139:40]
  assign io_actor_0_out_bits_write = block_blocked & block_blocked_1 ? _GEN_200 : io_actor_0_in_bits_write; // @[LockPool.scala 139:40]
  assign io_actor_0_out_bits_address = block_blocked & block_blocked_1 ? _GEN_202 : io_actor_0_in_bits_address; // @[LockPool.scala 139:40]
  assign io_actor_0_out_bits_size = block_blocked & block_blocked_1 ? _GEN_204 : io_actor_0_in_bits_size; // @[LockPool.scala 139:40]
  assign io_actor_0_out_bits_stride = block_blocked & block_blocked_1 ? _GEN_206 : io_actor_0_in_bits_stride; // @[LockPool.scala 139:40]
  assign io_actor_0_out_bits_reverse = block_blocked & block_blocked_1 ? _GEN_208 : io_actor_0_in_bits_reverse; // @[LockPool.scala 139:40]
  assign io_actor_1_in_ready = block_blocked & block_blocked_1 ? _GEN_195 : _GEN_15; // @[LockPool.scala 139:40]
  assign io_actor_1_out_valid = block_blocked & block_blocked_1 ? _GEN_199 : _GEN_16; // @[LockPool.scala 139:40]
  assign io_actor_1_out_bits_write = block_blocked & block_blocked_1 ? _GEN_201 : io_actor_1_in_bits_write; // @[LockPool.scala 139:40]
  assign io_actor_1_out_bits_address = block_blocked & block_blocked_1 ? _GEN_203 : io_actor_1_in_bits_address; // @[LockPool.scala 139:40]
  assign io_actor_1_out_bits_size = block_blocked & block_blocked_1 ? _GEN_205 : io_actor_1_in_bits_size; // @[LockPool.scala 139:40]
  assign io_actor_1_out_bits_stride = block_blocked & block_blocked_1 ? _GEN_207 : io_actor_1_in_bits_stride; // @[LockPool.scala 139:40]
  assign io_actor_1_out_bits_reverse = block_blocked & block_blocked_1 & _GEN_209; // @[LockPool.scala 139:40]
  assign io_lock_ready = ~(_GEN_39 & io_lock_bits_by != _GEN_37); // @[LockPool.scala 104:24]
  always @(posedge clock) begin
    if (reset) begin // @[LockPool.scala 55:21]
      lock_0_cond_write <= 1'h0; // @[LockPool.scala 55:21]
    end else if (lock_0_held) begin // @[LockPool.scala 108:18]
      if (observed) begin // @[LockPool.scala 109:22]
        if (incoming) begin // @[LockPool.scala 110:24]
          lock_0_cond_write <= _GEN_63;
        end
      end else if (incoming) begin // @[LockPool.scala 122:24]
        lock_0_cond_write <= _GEN_78;
      end
    end else if (incoming) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_0_cond_write <= _GEN_56;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_0_cond_address <= 14'h0; // @[LockPool.scala 55:21]
    end else if (lock_0_held) begin // @[LockPool.scala 108:18]
      if (observed) begin // @[LockPool.scala 109:22]
        if (incoming) begin // @[LockPool.scala 110:24]
          lock_0_cond_address <= _GEN_64;
        end
      end else if (incoming) begin // @[LockPool.scala 122:24]
        lock_0_cond_address <= _GEN_79;
      end
    end else if (incoming) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_0_cond_address <= _GEN_57;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_0_cond_size <= 14'h0; // @[LockPool.scala 55:21]
    end else if (lock_0_held) begin // @[LockPool.scala 108:18]
      if (observed) begin // @[LockPool.scala 109:22]
        if (incoming) begin // @[LockPool.scala 110:24]
          lock_0_cond_size <= _GEN_65;
        end
      end else if (incoming) begin // @[LockPool.scala 122:24]
        lock_0_cond_size <= _GEN_80;
      end
    end else if (incoming) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_0_cond_size <= _GEN_58;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_0_cond_stride <= 3'h0; // @[LockPool.scala 55:21]
    end else if (lock_0_held) begin // @[LockPool.scala 108:18]
      if (observed) begin // @[LockPool.scala 109:22]
        if (incoming) begin // @[LockPool.scala 110:24]
          lock_0_cond_stride <= _GEN_66;
        end
      end else if (incoming) begin // @[LockPool.scala 122:24]
        lock_0_cond_stride <= _GEN_81;
      end
    end else if (incoming) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_0_cond_stride <= _GEN_59;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_0_cond_reverse <= 1'h0; // @[LockPool.scala 55:21]
    end else if (lock_0_held) begin // @[LockPool.scala 108:18]
      if (observed) begin // @[LockPool.scala 109:22]
        if (incoming) begin // @[LockPool.scala 110:24]
          lock_0_cond_reverse <= _GEN_67;
        end
      end else if (incoming) begin // @[LockPool.scala 122:24]
        lock_0_cond_reverse <= _GEN_82;
      end
    end else if (incoming) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_0_cond_reverse <= _GEN_60;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_0_held <= 1'h0; // @[LockPool.scala 55:21]
    end else if (lock_0_held) begin // @[LockPool.scala 108:18]
      if (observed) begin // @[LockPool.scala 109:22]
        lock_0_held <= _GEN_68;
      end else if (incoming) begin // @[LockPool.scala 122:24]
        lock_0_held <= _GEN_76;
      end
    end else if (incoming) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_0_held <= _GEN_75;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_0_by <= 1'h0; // @[LockPool.scala 55:21]
    end else if (lock_0_held) begin // @[LockPool.scala 108:18]
      if (observed) begin // @[LockPool.scala 109:22]
        if (incoming) begin // @[LockPool.scala 110:24]
          lock_0_by <= _GEN_62;
        end
      end else if (incoming) begin // @[LockPool.scala 122:24]
        lock_0_by <= _GEN_77;
      end
    end else if (incoming) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_0_by <= _GEN_55;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_1_cond_write <= 1'h0; // @[LockPool.scala 55:21]
    end else if (lock_1_held) begin // @[LockPool.scala 108:18]
      if (observed_1) begin // @[LockPool.scala 109:22]
        if (io_lock_bits_lock) begin // @[LockPool.scala 110:24]
          lock_1_cond_write <= _GEN_139;
        end
      end else if (io_lock_bits_lock) begin // @[LockPool.scala 122:24]
        lock_1_cond_write <= _GEN_154;
      end
    end else if (io_lock_bits_lock) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_1_cond_write <= _GEN_133;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_1_cond_address <= 14'h0; // @[LockPool.scala 55:21]
    end else if (lock_1_held) begin // @[LockPool.scala 108:18]
      if (observed_1) begin // @[LockPool.scala 109:22]
        if (io_lock_bits_lock) begin // @[LockPool.scala 110:24]
          lock_1_cond_address <= _GEN_140;
        end
      end else if (io_lock_bits_lock) begin // @[LockPool.scala 122:24]
        lock_1_cond_address <= _GEN_155;
      end
    end else if (io_lock_bits_lock) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_1_cond_address <= _GEN_134;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_1_cond_size <= 14'h0; // @[LockPool.scala 55:21]
    end else if (lock_1_held) begin // @[LockPool.scala 108:18]
      if (observed_1) begin // @[LockPool.scala 109:22]
        if (io_lock_bits_lock) begin // @[LockPool.scala 110:24]
          lock_1_cond_size <= _GEN_141;
        end
      end else if (io_lock_bits_lock) begin // @[LockPool.scala 122:24]
        lock_1_cond_size <= _GEN_156;
      end
    end else if (io_lock_bits_lock) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_1_cond_size <= _GEN_135;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_1_cond_stride <= 3'h0; // @[LockPool.scala 55:21]
    end else if (lock_1_held) begin // @[LockPool.scala 108:18]
      if (observed_1) begin // @[LockPool.scala 109:22]
        if (io_lock_bits_lock) begin // @[LockPool.scala 110:24]
          lock_1_cond_stride <= _GEN_142;
        end
      end else if (io_lock_bits_lock) begin // @[LockPool.scala 122:24]
        lock_1_cond_stride <= _GEN_157;
      end
    end else if (io_lock_bits_lock) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_1_cond_stride <= _GEN_136;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_1_cond_reverse <= 1'h0; // @[LockPool.scala 55:21]
    end else if (lock_1_held) begin // @[LockPool.scala 108:18]
      if (observed_1) begin // @[LockPool.scala 109:22]
        if (io_lock_bits_lock) begin // @[LockPool.scala 110:24]
          lock_1_cond_reverse <= _GEN_143;
        end
      end else if (io_lock_bits_lock) begin // @[LockPool.scala 122:24]
        lock_1_cond_reverse <= _GEN_158;
      end
    end else if (io_lock_bits_lock) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_1_cond_reverse <= _GEN_137;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_1_held <= 1'h0; // @[LockPool.scala 55:21]
    end else if (lock_1_held) begin // @[LockPool.scala 108:18]
      if (observed_1) begin // @[LockPool.scala 109:22]
        lock_1_held <= _GEN_144;
      end else if (io_lock_bits_lock) begin // @[LockPool.scala 122:24]
        lock_1_held <= _GEN_152;
      end
    end else if (io_lock_bits_lock) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_1_held <= _GEN_151;
      end
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_1_by <= 1'h0; // @[LockPool.scala 55:21]
    end else if (lock_1_held) begin // @[LockPool.scala 108:18]
      if (observed_1) begin // @[LockPool.scala 109:22]
        if (io_lock_bits_lock) begin // @[LockPool.scala 110:24]
          lock_1_by <= _GEN_138;
        end
      end else if (io_lock_bits_lock) begin // @[LockPool.scala 122:24]
        lock_1_by <= _GEN_153;
      end
    end else if (io_lock_bits_lock) begin // @[LockPool.scala 130:22]
      if (~incomingObserved) begin // @[LockPool.scala 131:33]
        lock_1_by <= _GEN_132;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lock_0_cond_write = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  lock_0_cond_address = _RAND_1[13:0];
  _RAND_2 = {1{`RANDOM}};
  lock_0_cond_size = _RAND_2[13:0];
  _RAND_3 = {1{`RANDOM}};
  lock_0_cond_stride = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  lock_0_cond_reverse = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lock_0_held = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lock_0_by = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lock_1_cond_write = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  lock_1_cond_address = _RAND_8[13:0];
  _RAND_9 = {1{`RANDOM}};
  lock_1_cond_size = _RAND_9[13:0];
  _RAND_10 = {1{`RANDOM}};
  lock_1_cond_stride = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  lock_1_cond_reverse = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lock_1_held = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lock_1_by = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Counter_4(
  input         clock,
  input         reset,
  input         io_value_ready,
  output [11:0] io_value_bits,
  input         io_resetValue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [11:0] value; // @[Counter.scala 16:22]
  wire [11:0] _value_T_1 = value + 12'h1; // @[Counter.scala 24:22]
  assign io_value_bits = value; // @[Counter.scala 18:17]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 16:22]
      value <= 12'h0; // @[Counter.scala 16:22]
    end else if (io_resetValue) begin // @[Counter.scala 27:23]
      value <= 12'h0; // @[Counter.scala 28:11]
    end else if (io_value_ready) begin // @[Counter.scala 20:24]
      if (value == 12'hfff) begin // @[Counter.scala 21:31]
        value <= 12'h0; // @[Counter.scala 22:13]
      end else begin
        value <= _value_T_1; // @[Counter.scala 24:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CountBy_4(
  input         clock,
  input         reset,
  input         io_value_ready,
  output [11:0] io_value_bits,
  input  [11:0] io_step,
  input         io_resetValue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [11:0] value; // @[CountBy.scala 17:22]
  wire [12:0] _GEN_3 = {{1'd0}, io_step}; // @[CountBy.scala 22:24]
  wire [12:0] _T_1 = 13'h1000 - _GEN_3; // @[CountBy.scala 22:24]
  wire [12:0] _GEN_4 = {{1'd0}, value}; // @[CountBy.scala 22:16]
  wire [11:0] _value_T_1 = value + io_step; // @[CountBy.scala 25:22]
  assign io_value_bits = value; // @[CountBy.scala 19:17]
  always @(posedge clock) begin
    if (reset) begin // @[CountBy.scala 17:22]
      value <= 12'h0; // @[CountBy.scala 17:22]
    end else if (io_resetValue) begin // @[CountBy.scala 28:23]
      value <= 12'h0; // @[CountBy.scala 29:11]
    end else if (io_value_ready) begin // @[CountBy.scala 21:24]
      if (_GEN_4 >= _T_1) begin // @[CountBy.scala 22:36]
        value <= 12'h0; // @[CountBy.scala 23:13]
      end else begin
        value <= _value_T_1; // @[CountBy.scala 25:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SizeAndStrideHandler_4(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [3:0]  io_in_bits_instruction_op,
  input         io_in_bits_instruction_sourceLeft,
  input         io_in_bits_instruction_sourceRight,
  input         io_in_bits_instruction_dest,
  input  [11:0] io_in_bits_address,
  input  [11:0] io_in_bits_altAddress,
  input         io_in_bits_read,
  input         io_in_bits_write,
  input         io_in_bits_accumulate,
  input  [11:0] io_in_bits_size,
  input  [2:0]  io_in_bits_stride,
  input         io_in_bits_reverse,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_instruction_op,
  output        io_out_bits_instruction_sourceLeft,
  output        io_out_bits_instruction_sourceRight,
  output        io_out_bits_instruction_dest,
  output [11:0] io_out_bits_address,
  output [11:0] io_out_bits_altAddress,
  output        io_out_bits_read,
  output        io_out_bits_write,
  output        io_out_bits_accumulate
);
  wire  sizeCounter_clock; // @[Counter.scala 34:19]
  wire  sizeCounter_reset; // @[Counter.scala 34:19]
  wire  sizeCounter_io_value_ready; // @[Counter.scala 34:19]
  wire [11:0] sizeCounter_io_value_bits; // @[Counter.scala 34:19]
  wire  sizeCounter_io_resetValue; // @[Counter.scala 34:19]
  wire  addressCounter_clock; // @[CountBy.scala 35:19]
  wire  addressCounter_reset; // @[CountBy.scala 35:19]
  wire  addressCounter_io_value_ready; // @[CountBy.scala 35:19]
  wire [11:0] addressCounter_io_value_bits; // @[CountBy.scala 35:19]
  wire [11:0] addressCounter_io_step; // @[CountBy.scala 35:19]
  wire  addressCounter_io_resetValue; // @[CountBy.scala 35:19]
  wire [7:0] stride = 8'h1 << io_in_bits_stride; // @[SizeAndStrideHandler.scala 30:20]
  wire [11:0] _io_out_bits_address_T_1 = io_in_bits_address - addressCounter_io_value_bits; // @[SizeAndStrideHandler.scala 46:44]
  wire [11:0] _io_out_bits_address_T_3 = io_in_bits_address + addressCounter_io_value_bits; // @[SizeAndStrideHandler.scala 48:44]
  wire  fire = io_in_valid & io_out_ready; // @[SizeAndStrideHandler.scala 51:23]
  Counter_4 sizeCounter ( // @[Counter.scala 34:19]
    .clock(sizeCounter_clock),
    .reset(sizeCounter_reset),
    .io_value_ready(sizeCounter_io_value_ready),
    .io_value_bits(sizeCounter_io_value_bits),
    .io_resetValue(sizeCounter_io_resetValue)
  );
  CountBy_4 addressCounter ( // @[CountBy.scala 35:19]
    .clock(addressCounter_clock),
    .reset(addressCounter_reset),
    .io_value_ready(addressCounter_io_value_ready),
    .io_value_bits(addressCounter_io_value_bits),
    .io_step(addressCounter_io_step),
    .io_resetValue(addressCounter_io_resetValue)
  );
  assign io_in_ready = sizeCounter_io_value_bits == io_in_bits_size & io_out_ready; // @[SizeAndStrideHandler.scala 53:52 54:14 58:14]
  assign io_out_valid = io_in_valid; // @[SizeAndStrideHandler.scala 35:16]
  assign io_out_bits_instruction_op = io_in_bits_instruction_op; // @[SizeAndStrideHandler.scala 38:34]
  assign io_out_bits_instruction_sourceLeft = io_in_bits_instruction_sourceLeft; // @[SizeAndStrideHandler.scala 38:34]
  assign io_out_bits_instruction_sourceRight = io_in_bits_instruction_sourceRight; // @[SizeAndStrideHandler.scala 38:34]
  assign io_out_bits_instruction_dest = io_in_bits_instruction_dest; // @[SizeAndStrideHandler.scala 38:34]
  assign io_out_bits_address = io_in_bits_reverse ? _io_out_bits_address_T_1 : _io_out_bits_address_T_3; // @[SizeAndStrideHandler.scala 45:25 46:25 48:25]
  assign io_out_bits_altAddress = io_in_bits_altAddress; // @[SizeAndStrideHandler.scala 38:34]
  assign io_out_bits_read = io_in_bits_read; // @[SizeAndStrideHandler.scala 38:34]
  assign io_out_bits_write = io_in_bits_write; // @[SizeAndStrideHandler.scala 38:34]
  assign io_out_bits_accumulate = io_in_bits_accumulate; // @[SizeAndStrideHandler.scala 38:34]
  assign sizeCounter_clock = clock;
  assign sizeCounter_reset = reset;
  assign sizeCounter_io_value_ready = sizeCounter_io_value_bits == io_in_bits_size ? 1'h0 : fire; // @[Counter.scala 36:22 SizeAndStrideHandler.scala 53:52 59:32]
  assign sizeCounter_io_resetValue = sizeCounter_io_value_bits == io_in_bits_size & fire; // @[Counter.scala 35:21 SizeAndStrideHandler.scala 53:52 55:31]
  assign addressCounter_clock = clock;
  assign addressCounter_reset = reset;
  assign addressCounter_io_value_ready = sizeCounter_io_value_bits == io_in_bits_size ? 1'h0 : fire; // @[Counter.scala 36:22 SizeAndStrideHandler.scala 53:52 59:32]
  assign addressCounter_io_step = {{4'd0}, stride}; // @[CountBy.scala 36:15]
  assign addressCounter_io_resetValue = sizeCounter_io_value_bits == io_in_bits_size & fire; // @[Counter.scala 35:21 SizeAndStrideHandler.scala 53:52 55:31]
endmodule
module Queue_4(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_instruction_op,
  input         io_enq_bits_instruction_sourceLeft,
  input         io_enq_bits_instruction_sourceRight,
  input         io_enq_bits_instruction_dest,
  input  [11:0] io_enq_bits_address,
  input  [11:0] io_enq_bits_altAddress,
  input         io_enq_bits_read,
  input         io_enq_bits_write,
  input         io_enq_bits_accumulate,
  input  [11:0] io_enq_bits_size,
  input  [2:0]  io_enq_bits_stride,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_instruction_op,
  output        io_deq_bits_instruction_sourceLeft,
  output        io_deq_bits_instruction_sourceRight,
  output        io_deq_bits_instruction_dest,
  output [11:0] io_deq_bits_address,
  output [11:0] io_deq_bits_altAddress,
  output        io_deq_bits_read,
  output        io_deq_bits_write,
  output        io_deq_bits_accumulate,
  output [11:0] io_deq_bits_size,
  output [2:0]  io_deq_bits_stride,
  output        io_deq_bits_reverse
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_instruction_op [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_instruction_op_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_instruction_op_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_instruction_op_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_instruction_op_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_instruction_op_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_op_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_instruction_op_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_instruction_sourceLeft [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_instruction_sourceLeft_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_instruction_sourceLeft_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_instruction_sourceRight [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_instruction_sourceRight_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_instruction_sourceRight_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_instruction_dest [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_instruction_dest_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_instruction_dest_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_MPORT_en; // @[Decoupled.scala 259:95]
  reg [11:0] ram_address [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [11:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [11:0] ram_address_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_address_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 259:95]
  reg [11:0] ram_altAddress [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_altAddress_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_altAddress_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [11:0] ram_altAddress_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [11:0] ram_altAddress_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_altAddress_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_altAddress_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_altAddress_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_read [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_read_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_read_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_read_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_read_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_write [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_write_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_write_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_accumulate [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_accumulate_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_accumulate_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_MPORT_en; // @[Decoupled.scala 259:95]
  reg [11:0] ram_size [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [11:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [11:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_stride [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_stride_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_stride_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_stride_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_stride_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_stride_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_stride_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_stride_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_reverse [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_reverse_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_reverse_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_reverse_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_reverse_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_reverse_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_reverse_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_reverse_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [5:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [5:0] _value_T_1 = enq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire  _GEN_23 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_23 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire [5:0] _value_T_3 = deq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_instruction_op_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instruction_op_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instruction_op_io_deq_bits_MPORT_data = ram_instruction_op[ram_instruction_op_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_instruction_op_MPORT_data = io_enq_bits_instruction_op;
  assign ram_instruction_op_MPORT_addr = enq_ptr_value;
  assign ram_instruction_op_MPORT_mask = 1'h1;
  assign ram_instruction_op_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_instruction_sourceLeft_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instruction_sourceLeft_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instruction_sourceLeft_io_deq_bits_MPORT_data =
    ram_instruction_sourceLeft[ram_instruction_sourceLeft_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_instruction_sourceLeft_MPORT_data = io_enq_bits_instruction_sourceLeft;
  assign ram_instruction_sourceLeft_MPORT_addr = enq_ptr_value;
  assign ram_instruction_sourceLeft_MPORT_mask = 1'h1;
  assign ram_instruction_sourceLeft_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_instruction_sourceRight_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instruction_sourceRight_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instruction_sourceRight_io_deq_bits_MPORT_data =
    ram_instruction_sourceRight[ram_instruction_sourceRight_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_instruction_sourceRight_MPORT_data = io_enq_bits_instruction_sourceRight;
  assign ram_instruction_sourceRight_MPORT_addr = enq_ptr_value;
  assign ram_instruction_sourceRight_MPORT_mask = 1'h1;
  assign ram_instruction_sourceRight_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_instruction_dest_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instruction_dest_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instruction_dest_io_deq_bits_MPORT_data = ram_instruction_dest[ram_instruction_dest_io_deq_bits_MPORT_addr]
    ; // @[Decoupled.scala 259:95]
  assign ram_instruction_dest_MPORT_data = io_enq_bits_instruction_dest;
  assign ram_instruction_dest_MPORT_addr = enq_ptr_value;
  assign ram_instruction_dest_MPORT_mask = 1'h1;
  assign ram_instruction_dest_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = enq_ptr_value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_altAddress_io_deq_bits_MPORT_en = 1'h1;
  assign ram_altAddress_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_altAddress_io_deq_bits_MPORT_data = ram_altAddress[ram_altAddress_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_altAddress_MPORT_data = io_enq_bits_altAddress;
  assign ram_altAddress_MPORT_addr = enq_ptr_value;
  assign ram_altAddress_MPORT_mask = 1'h1;
  assign ram_altAddress_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_read_io_deq_bits_MPORT_en = 1'h1;
  assign ram_read_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_read_io_deq_bits_MPORT_data = ram_read[ram_read_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_read_MPORT_data = io_enq_bits_read;
  assign ram_read_MPORT_addr = enq_ptr_value;
  assign ram_read_MPORT_mask = 1'h1;
  assign ram_read_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_write_io_deq_bits_MPORT_en = 1'h1;
  assign ram_write_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_write_io_deq_bits_MPORT_data = ram_write[ram_write_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_write_MPORT_data = io_enq_bits_write;
  assign ram_write_MPORT_addr = enq_ptr_value;
  assign ram_write_MPORT_mask = 1'h1;
  assign ram_write_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_accumulate_io_deq_bits_MPORT_en = 1'h1;
  assign ram_accumulate_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_accumulate_io_deq_bits_MPORT_data = ram_accumulate[ram_accumulate_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_accumulate_MPORT_data = io_enq_bits_accumulate;
  assign ram_accumulate_MPORT_addr = enq_ptr_value;
  assign ram_accumulate_MPORT_mask = 1'h1;
  assign ram_accumulate_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_stride_io_deq_bits_MPORT_en = 1'h1;
  assign ram_stride_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_stride_io_deq_bits_MPORT_data = ram_stride[ram_stride_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_stride_MPORT_data = io_enq_bits_stride;
  assign ram_stride_MPORT_addr = enq_ptr_value;
  assign ram_stride_MPORT_mask = 1'h1;
  assign ram_stride_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_reverse_io_deq_bits_MPORT_en = 1'h1;
  assign ram_reverse_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_reverse_io_deq_bits_MPORT_data = ram_reverse[ram_reverse_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_reverse_MPORT_data = 1'h0;
  assign ram_reverse_MPORT_addr = enq_ptr_value;
  assign ram_reverse_MPORT_mask = 1'h1;
  assign ram_reverse_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | ~full; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_instruction_op = empty ? io_enq_bits_instruction_op : ram_instruction_op_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_instruction_sourceLeft = empty ? io_enq_bits_instruction_sourceLeft :
    ram_instruction_sourceLeft_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_instruction_sourceRight = empty ? io_enq_bits_instruction_sourceRight :
    ram_instruction_sourceRight_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_instruction_dest = empty ? io_enq_bits_instruction_dest :
    ram_instruction_dest_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_address = empty ? io_enq_bits_address : ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_altAddress = empty ? io_enq_bits_altAddress : ram_altAddress_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_read = empty ? io_enq_bits_read : ram_read_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_write = empty ? io_enq_bits_write : ram_write_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_accumulate = empty ? io_enq_bits_accumulate : ram_accumulate_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_stride = empty ? io_enq_bits_stride : ram_stride_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_reverse = empty ? 1'h0 : ram_reverse_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_instruction_op_MPORT_en & ram_instruction_op_MPORT_mask) begin
      ram_instruction_op[ram_instruction_op_MPORT_addr] <= ram_instruction_op_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_instruction_sourceLeft_MPORT_en & ram_instruction_sourceLeft_MPORT_mask) begin
      ram_instruction_sourceLeft[ram_instruction_sourceLeft_MPORT_addr] <= ram_instruction_sourceLeft_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_instruction_sourceRight_MPORT_en & ram_instruction_sourceRight_MPORT_mask) begin
      ram_instruction_sourceRight[ram_instruction_sourceRight_MPORT_addr] <= ram_instruction_sourceRight_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_instruction_dest_MPORT_en & ram_instruction_dest_MPORT_mask) begin
      ram_instruction_dest[ram_instruction_dest_MPORT_addr] <= ram_instruction_dest_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_altAddress_MPORT_en & ram_altAddress_MPORT_mask) begin
      ram_altAddress[ram_altAddress_MPORT_addr] <= ram_altAddress_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_read_MPORT_en & ram_read_MPORT_mask) begin
      ram_read[ram_read_MPORT_addr] <= ram_read_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_write_MPORT_en & ram_write_MPORT_mask) begin
      ram_write[ram_write_MPORT_addr] <= ram_write_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_accumulate_MPORT_en & ram_accumulate_MPORT_mask) begin
      ram_accumulate[ram_accumulate_MPORT_addr] <= ram_accumulate_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_stride_MPORT_en & ram_stride_MPORT_mask) begin
      ram_stride[ram_stride_MPORT_addr] <= ram_stride_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_reverse_MPORT_en & ram_reverse_MPORT_mask) begin
      ram_reverse[ram_reverse_MPORT_addr] <= ram_reverse_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_instruction_op[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_instruction_sourceLeft[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_instruction_sourceRight[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_instruction_dest[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[11:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_altAddress[initvar] = _RAND_5[11:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_read[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_write[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_accumulate[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_size[initvar] = _RAND_9[11:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_stride[initvar] = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_reverse[initvar] = _RAND_11[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  enq_ptr_value = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  deq_ptr_value = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  maybe_full = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SizeHandler(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_load,
  input         io_in_bits_zeroes,
  input  [13:0] io_in_bits_size,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_load,
  output        io_out_bits_zeroes
);
  wire  sizeCounter_clock; // @[Counter.scala 34:19]
  wire  sizeCounter_reset; // @[Counter.scala 34:19]
  wire  sizeCounter_io_value_ready; // @[Counter.scala 34:19]
  wire [13:0] sizeCounter_io_value_bits; // @[Counter.scala 34:19]
  wire  sizeCounter_io_resetValue; // @[Counter.scala 34:19]
  wire  fire = io_in_valid & io_out_ready; // @[SizeHandler.scala 32:23]
  Counter_2 sizeCounter ( // @[Counter.scala 34:19]
    .clock(sizeCounter_clock),
    .reset(sizeCounter_reset),
    .io_value_ready(sizeCounter_io_value_ready),
    .io_value_bits(sizeCounter_io_value_bits),
    .io_resetValue(sizeCounter_io_resetValue)
  );
  assign io_in_ready = sizeCounter_io_value_bits == io_in_bits_size & io_out_ready; // @[SizeHandler.scala 34:52 35:14 38:14]
  assign io_out_valid = io_in_valid; // @[SizeHandler.scala 25:16]
  assign io_out_bits_load = io_in_bits_load; // @[SizeHandler.scala 28:34]
  assign io_out_bits_zeroes = io_in_bits_zeroes; // @[SizeHandler.scala 28:34]
  assign sizeCounter_clock = clock;
  assign sizeCounter_reset = reset;
  assign sizeCounter_io_value_ready = sizeCounter_io_value_bits == io_in_bits_size ? 1'h0 : fire; // @[SizeHandler.scala 34:52 Counter.scala 36:22 SizeHandler.scala 39:32]
  assign sizeCounter_io_resetValue = sizeCounter_io_value_bits == io_in_bits_size & fire; // @[SizeHandler.scala 34:52 Counter.scala 35:21 SizeHandler.scala 36:31]
endmodule
module Queue_5(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_load,
  input         io_enq_bits_zeroes,
  input  [13:0] io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_load,
  output        io_deq_bits_zeroes,
  output [13:0] io_deq_bits_size
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  ram_load [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_load_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_load_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_load_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_load_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_load_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_load_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_load_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_zeroes [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_zeroes_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_zeroes_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_MPORT_en; // @[Decoupled.scala 259:95]
  reg [13:0] ram_size [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [5:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [5:0] _value_T_1 = enq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire  _GEN_14 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_14 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire [5:0] _value_T_3 = deq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_load_io_deq_bits_MPORT_en = 1'h1;
  assign ram_load_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_load_io_deq_bits_MPORT_data = ram_load[ram_load_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_load_MPORT_data = io_enq_bits_load;
  assign ram_load_MPORT_addr = enq_ptr_value;
  assign ram_load_MPORT_mask = 1'h1;
  assign ram_load_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_zeroes_io_deq_bits_MPORT_en = 1'h1;
  assign ram_zeroes_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_zeroes_io_deq_bits_MPORT_data = ram_zeroes[ram_zeroes_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_zeroes_MPORT_data = io_enq_bits_zeroes;
  assign ram_zeroes_MPORT_addr = enq_ptr_value;
  assign ram_zeroes_MPORT_mask = 1'h1;
  assign ram_zeroes_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | ~full; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_load = empty ? io_enq_bits_load : ram_load_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_zeroes = empty ? io_enq_bits_zeroes : ram_zeroes_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_load_MPORT_en & ram_load_MPORT_mask) begin
      ram_load[ram_load_MPORT_addr] <= ram_load_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_zeroes_MPORT_en & ram_zeroes_MPORT_mask) begin
      ram_zeroes[ram_zeroes_MPORT_addr] <= ram_zeroes_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_load[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_zeroes[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[13:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_6(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_kind,
  input  [13:0] io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_kind,
  output [13:0] io_deq_bits_size
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_kind [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_kind_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_kind_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_kind_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_kind_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_kind_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_kind_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_kind_MPORT_en; // @[Decoupled.scala 259:95]
  reg [13:0] ram_size [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [5:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [5:0] _value_T_1 = enq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire  _GEN_13 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_13 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire [5:0] _value_T_3 = deq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_kind_io_deq_bits_MPORT_en = 1'h1;
  assign ram_kind_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_kind_io_deq_bits_MPORT_data = ram_kind[ram_kind_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_kind_MPORT_data = io_enq_bits_kind;
  assign ram_kind_MPORT_addr = enq_ptr_value;
  assign ram_kind_MPORT_mask = 1'h1;
  assign ram_kind_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | ~full; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_kind = empty ? io_enq_bits_kind : ram_kind_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_kind_MPORT_en & ram_kind_MPORT_mask) begin
      ram_kind[ram_kind_MPORT_addr] <= ram_kind_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_kind[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[13:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SizeHandler_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [1:0]  io_in_bits_kind,
  input  [13:0] io_in_bits_size,
  input         io_out_ready,
  output        io_out_valid,
  output [1:0]  io_out_bits_kind
);
  wire  sizeCounter_clock; // @[Counter.scala 34:19]
  wire  sizeCounter_reset; // @[Counter.scala 34:19]
  wire  sizeCounter_io_value_ready; // @[Counter.scala 34:19]
  wire [13:0] sizeCounter_io_value_bits; // @[Counter.scala 34:19]
  wire  sizeCounter_io_resetValue; // @[Counter.scala 34:19]
  wire  fire = io_in_valid & io_out_ready; // @[SizeHandler.scala 32:23]
  Counter_2 sizeCounter ( // @[Counter.scala 34:19]
    .clock(sizeCounter_clock),
    .reset(sizeCounter_reset),
    .io_value_ready(sizeCounter_io_value_ready),
    .io_value_bits(sizeCounter_io_value_bits),
    .io_resetValue(sizeCounter_io_resetValue)
  );
  assign io_in_ready = sizeCounter_io_value_bits == io_in_bits_size & io_out_ready; // @[SizeHandler.scala 34:52 35:14 38:14]
  assign io_out_valid = io_in_valid; // @[SizeHandler.scala 25:16]
  assign io_out_bits_kind = io_in_bits_kind; // @[SizeHandler.scala 28:34]
  assign sizeCounter_clock = clock;
  assign sizeCounter_reset = reset;
  assign sizeCounter_io_value_ready = sizeCounter_io_value_bits == io_in_bits_size ? 1'h0 : fire; // @[SizeHandler.scala 34:52 Counter.scala 36:22 SizeHandler.scala 39:32]
  assign sizeCounter_io_resetValue = sizeCounter_io_value_bits == io_in_bits_size & fire; // @[SizeHandler.scala 34:52 Counter.scala 35:21 SizeHandler.scala 36:31]
endmodule
module Queue_7(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_kind,
  input  [13:0] io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_kind,
  output [13:0] io_deq_bits_size
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_kind [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_kind_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_kind_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_kind_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_kind_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_kind_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_kind_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_kind_MPORT_en; // @[Decoupled.scala 259:95]
  reg [13:0] ram_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_10 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_10 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_kind_io_deq_bits_MPORT_en = 1'h1;
  assign ram_kind_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_kind_io_deq_bits_MPORT_data = ram_kind[ram_kind_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_kind_MPORT_data = io_enq_bits_kind;
  assign ram_kind_MPORT_addr = 1'h0;
  assign ram_kind_MPORT_mask = 1'h1;
  assign ram_kind_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_kind = empty ? io_enq_bits_kind : ram_kind_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_kind_MPORT_en & ram_kind_MPORT_mask) begin
      ram_kind[ram_kind_MPORT_addr] <= ram_kind_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_kind[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[13:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MultiEnqueue(
  input   clock,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input   io_out_0_ready,
  output  io_out_0_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  enq_0; // @[MultiEnqueue.scala 16:47]
  wire  allEnqueued = io_out_0_ready | enq_0; // @[MultiEnqueue.scala 22:34]
  wire  _io_out_0_valid_T = ~enq_0; // @[MultiEnqueue.scala 27:39]
  assign io_in_ready = io_out_0_ready | enq_0; // @[MultiEnqueue.scala 22:34]
  assign io_out_0_valid = io_in_valid & ~enq_0; // @[MultiEnqueue.scala 27:36]
  always @(posedge clock) begin
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_0 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_0 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_0_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_0 <= io_out_0_valid & io_out_0_ready; // @[MultiEnqueue.scala 32:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enq_0 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MultiEnqueue_1(
  input   clock,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input   io_out_0_ready,
  output  io_out_0_valid,
  input   io_out_1_ready,
  output  io_out_1_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  enq_0; // @[MultiEnqueue.scala 16:47]
  reg  enq_1; // @[MultiEnqueue.scala 16:47]
  wire  _allEnqueued_T = io_out_0_ready | enq_0; // @[MultiEnqueue.scala 22:34]
  wire  _allEnqueued_T_1 = io_out_1_ready | enq_1; // @[MultiEnqueue.scala 22:34]
  wire  allEnqueued = _allEnqueued_T & _allEnqueued_T_1; // @[MultiEnqueue.scala 24:15]
  wire  _io_out_0_valid_T = ~enq_0; // @[MultiEnqueue.scala 27:39]
  wire  _io_out_1_valid_T = ~enq_1; // @[MultiEnqueue.scala 27:39]
  assign io_in_ready = _allEnqueued_T & _allEnqueued_T_1; // @[MultiEnqueue.scala 24:15]
  assign io_out_0_valid = io_in_valid & ~enq_0; // @[MultiEnqueue.scala 27:36]
  assign io_out_1_valid = io_in_valid & ~enq_1; // @[MultiEnqueue.scala 27:36]
  always @(posedge clock) begin
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_0 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_0 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_0_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_0 <= io_out_0_valid & io_out_0_ready; // @[MultiEnqueue.scala 32:16]
    end
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_1 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_1 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_1_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_1 <= io_out_1_valid & io_out_1_ready; // @[MultiEnqueue.scala 32:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enq_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  enq_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MultiEnqueue_2(
  input   clock,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input   io_out_0_ready,
  output  io_out_0_valid,
  input   io_out_1_ready,
  output  io_out_1_valid,
  input   io_out_2_ready,
  output  io_out_2_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  enq_0; // @[MultiEnqueue.scala 16:47]
  reg  enq_1; // @[MultiEnqueue.scala 16:47]
  reg  enq_2; // @[MultiEnqueue.scala 16:47]
  wire  _allEnqueued_T = io_out_0_ready | enq_0; // @[MultiEnqueue.scala 22:34]
  wire  _allEnqueued_T_1 = io_out_1_ready | enq_1; // @[MultiEnqueue.scala 22:34]
  wire  _allEnqueued_T_2 = io_out_2_ready | enq_2; // @[MultiEnqueue.scala 22:34]
  wire  allEnqueued = _allEnqueued_T & _allEnqueued_T_1 & _allEnqueued_T_2; // @[MultiEnqueue.scala 24:15]
  wire  _io_out_0_valid_T = ~enq_0; // @[MultiEnqueue.scala 27:39]
  wire  _io_out_1_valid_T = ~enq_1; // @[MultiEnqueue.scala 27:39]
  wire  _io_out_2_valid_T = ~enq_2; // @[MultiEnqueue.scala 27:39]
  assign io_in_ready = _allEnqueued_T & _allEnqueued_T_1 & _allEnqueued_T_2; // @[MultiEnqueue.scala 24:15]
  assign io_out_0_valid = io_in_valid & ~enq_0; // @[MultiEnqueue.scala 27:36]
  assign io_out_1_valid = io_in_valid & ~enq_1; // @[MultiEnqueue.scala 27:36]
  assign io_out_2_valid = io_in_valid & ~enq_2; // @[MultiEnqueue.scala 27:36]
  always @(posedge clock) begin
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_0 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_0 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_0_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_0 <= io_out_0_valid & io_out_0_ready; // @[MultiEnqueue.scala 32:16]
    end
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_1 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_1 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_1_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_1 <= io_out_1_valid & io_out_1_ready; // @[MultiEnqueue.scala 32:16]
    end
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_2 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_2 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_2_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_2 <= io_out_2_valid & io_out_2_ready; // @[MultiEnqueue.scala 32:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enq_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  enq_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enq_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MultiEnqueue_3(
  input   clock,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input   io_out_0_ready,
  output  io_out_0_valid,
  input   io_out_1_ready,
  output  io_out_1_valid,
  input   io_out_2_ready,
  output  io_out_2_valid,
  input   io_out_3_ready,
  output  io_out_3_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  enq_0; // @[MultiEnqueue.scala 16:47]
  reg  enq_1; // @[MultiEnqueue.scala 16:47]
  reg  enq_2; // @[MultiEnqueue.scala 16:47]
  reg  enq_3; // @[MultiEnqueue.scala 16:47]
  wire  _allEnqueued_T = io_out_0_ready | enq_0; // @[MultiEnqueue.scala 22:34]
  wire  _allEnqueued_T_1 = io_out_1_ready | enq_1; // @[MultiEnqueue.scala 22:34]
  wire  _allEnqueued_T_2 = io_out_2_ready | enq_2; // @[MultiEnqueue.scala 22:34]
  wire  _allEnqueued_T_3 = io_out_3_ready | enq_3; // @[MultiEnqueue.scala 22:34]
  wire  allEnqueued = _allEnqueued_T & _allEnqueued_T_1 & _allEnqueued_T_2 & _allEnqueued_T_3; // @[MultiEnqueue.scala 24:15]
  wire  _io_out_0_valid_T = ~enq_0; // @[MultiEnqueue.scala 27:39]
  wire  _io_out_1_valid_T = ~enq_1; // @[MultiEnqueue.scala 27:39]
  wire  _io_out_2_valid_T = ~enq_2; // @[MultiEnqueue.scala 27:39]
  wire  _io_out_3_valid_T = ~enq_3; // @[MultiEnqueue.scala 27:39]
  assign io_in_ready = _allEnqueued_T & _allEnqueued_T_1 & _allEnqueued_T_2 & _allEnqueued_T_3; // @[MultiEnqueue.scala 24:15]
  assign io_out_0_valid = io_in_valid & ~enq_0; // @[MultiEnqueue.scala 27:36]
  assign io_out_1_valid = io_in_valid & ~enq_1; // @[MultiEnqueue.scala 27:36]
  assign io_out_2_valid = io_in_valid & ~enq_2; // @[MultiEnqueue.scala 27:36]
  assign io_out_3_valid = io_in_valid & ~enq_3; // @[MultiEnqueue.scala 27:36]
  always @(posedge clock) begin
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_0 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_0 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_0_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_0 <= io_out_0_valid & io_out_0_ready; // @[MultiEnqueue.scala 32:16]
    end
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_1 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_1 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_1_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_1 <= io_out_1_valid & io_out_1_ready; // @[MultiEnqueue.scala 32:16]
    end
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_2 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_2 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_2_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_2 <= io_out_2_valid & io_out_2_ready; // @[MultiEnqueue.scala 32:16]
    end
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_3 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_3 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_3_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_3 <= io_out_3_valid & io_out_3_ready; // @[MultiEnqueue.scala 32:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enq_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  enq_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enq_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enq_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MultiEnqueue_4(
  input   clock,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input   io_out_0_ready,
  output  io_out_0_valid,
  input   io_out_1_ready,
  output  io_out_1_valid,
  input   io_out_2_ready,
  output  io_out_2_valid,
  input   io_out_3_ready,
  output  io_out_3_valid,
  input   io_out_4_ready,
  output  io_out_4_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  enq_0; // @[MultiEnqueue.scala 16:47]
  reg  enq_1; // @[MultiEnqueue.scala 16:47]
  reg  enq_2; // @[MultiEnqueue.scala 16:47]
  reg  enq_3; // @[MultiEnqueue.scala 16:47]
  reg  enq_4; // @[MultiEnqueue.scala 16:47]
  wire  _allEnqueued_T = io_out_0_ready | enq_0; // @[MultiEnqueue.scala 22:34]
  wire  _allEnqueued_T_1 = io_out_1_ready | enq_1; // @[MultiEnqueue.scala 22:34]
  wire  _allEnqueued_T_2 = io_out_2_ready | enq_2; // @[MultiEnqueue.scala 22:34]
  wire  _allEnqueued_T_3 = io_out_3_ready | enq_3; // @[MultiEnqueue.scala 22:34]
  wire  _allEnqueued_T_4 = io_out_4_ready | enq_4; // @[MultiEnqueue.scala 22:34]
  wire  allEnqueued = _allEnqueued_T & _allEnqueued_T_1 & _allEnqueued_T_2 & _allEnqueued_T_3 & _allEnqueued_T_4; // @[MultiEnqueue.scala 24:15]
  wire  _io_out_0_valid_T = ~enq_0; // @[MultiEnqueue.scala 27:39]
  wire  _io_out_1_valid_T = ~enq_1; // @[MultiEnqueue.scala 27:39]
  wire  _io_out_2_valid_T = ~enq_2; // @[MultiEnqueue.scala 27:39]
  wire  _io_out_3_valid_T = ~enq_3; // @[MultiEnqueue.scala 27:39]
  wire  _io_out_4_valid_T = ~enq_4; // @[MultiEnqueue.scala 27:39]
  assign io_in_ready = _allEnqueued_T & _allEnqueued_T_1 & _allEnqueued_T_2 & _allEnqueued_T_3 & _allEnqueued_T_4; // @[MultiEnqueue.scala 24:15]
  assign io_out_0_valid = io_in_valid & ~enq_0; // @[MultiEnqueue.scala 27:36]
  assign io_out_1_valid = io_in_valid & ~enq_1; // @[MultiEnqueue.scala 27:36]
  assign io_out_2_valid = io_in_valid & ~enq_2; // @[MultiEnqueue.scala 27:36]
  assign io_out_3_valid = io_in_valid & ~enq_3; // @[MultiEnqueue.scala 27:36]
  assign io_out_4_valid = io_in_valid & ~enq_4; // @[MultiEnqueue.scala 27:36]
  always @(posedge clock) begin
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_0 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_0 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_0_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_0 <= io_out_0_valid & io_out_0_ready; // @[MultiEnqueue.scala 32:16]
    end
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_1 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_1 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_1_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_1 <= io_out_1_valid & io_out_1_ready; // @[MultiEnqueue.scala 32:16]
    end
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_2 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_2 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_2_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_2 <= io_out_2_valid & io_out_2_ready; // @[MultiEnqueue.scala 32:16]
    end
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_3 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_3 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_3_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_3 <= io_out_3_valid & io_out_3_ready; // @[MultiEnqueue.scala 32:16]
    end
    if (reset) begin // @[MultiEnqueue.scala 16:47]
      enq_4 <= 1'h0; // @[MultiEnqueue.scala 16:47]
    end else if (allEnqueued) begin // @[MultiEnqueue.scala 28:23]
      enq_4 <= 1'h0; // @[MultiEnqueue.scala 29:14]
    end else if (_io_out_4_valid_T) begin // @[MultiEnqueue.scala 31:21]
      enq_4 <= io_out_4_valid & io_out_4_ready; // @[MultiEnqueue.scala 32:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enq_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  enq_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enq_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enq_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  enq_4 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decoder(
  input         clock,
  input         reset,
  output        io_instruction_ready,
  input         io_instruction_valid,
  input  [3:0]  io_instruction_bits_opcode,
  input  [3:0]  io_instruction_bits_flags,
  input  [63:0] io_instruction_bits_arguments,
  input         io_memPortA_ready,
  output        io_memPortA_valid,
  output        io_memPortA_bits_write,
  output [13:0] io_memPortA_bits_address,
  input         io_memPortB_ready,
  output        io_memPortB_valid,
  output        io_memPortB_bits_write,
  output [13:0] io_memPortB_bits_address,
  input         io_dram0_ready,
  output        io_dram0_valid,
  output        io_dram0_bits_write,
  output [20:0] io_dram0_bits_address,
  output [20:0] io_dram0_bits_size,
  input         io_dram1_ready,
  output        io_dram1_valid,
  output        io_dram1_bits_write,
  output [20:0] io_dram1_bits_address,
  output [20:0] io_dram1_bits_size,
  input         io_dataflow_ready,
  output        io_dataflow_valid,
  output [3:0]  io_dataflow_bits_kind,
  output [13:0] io_dataflow_bits_size,
  input         io_hostDataflow_ready,
  output        io_hostDataflow_valid,
  output [1:0]  io_hostDataflow_bits_kind,
  input         io_acc_ready,
  output        io_acc_valid,
  output [3:0]  io_acc_bits_instruction_op,
  output        io_acc_bits_instruction_sourceLeft,
  output        io_acc_bits_instruction_sourceRight,
  output        io_acc_bits_instruction_dest,
  output [11:0] io_acc_bits_readAddress,
  output [11:0] io_acc_bits_writeAddress,
  output        io_acc_bits_accumulate,
  output        io_acc_bits_write,
  output        io_acc_bits_read,
  input         io_array_ready,
  output        io_array_valid,
  output        io_array_bits_load,
  output        io_array_bits_zeroes,
  output [31:0] io_config_dram0AddressOffset,
  output [3:0]  io_config_dram0CacheBehaviour,
  output [31:0] io_config_dram1AddressOffset,
  output [3:0]  io_config_dram1CacheBehaviour,
  output        io_timeout,
  output        io_error,
  output        io_tracepoint,
  output [31:0] io_programCounter
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  instruction_clock; // @[Decoupled.scala 361:21]
  wire  instruction_reset; // @[Decoupled.scala 361:21]
  wire  instruction_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  instruction_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [3:0] instruction_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] instruction_io_enq_bits_flags; // @[Decoupled.scala 361:21]
  wire [63:0] instruction_io_enq_bits_arguments; // @[Decoupled.scala 361:21]
  wire  instruction_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  instruction_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [3:0] instruction_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] instruction_io_deq_bits_flags; // @[Decoupled.scala 361:21]
  wire [63:0] instruction_io_deq_bits_arguments; // @[Decoupled.scala 361:21]
  wire  dram0Handler_clock; // @[Decoder.scala 144:28]
  wire  dram0Handler_reset; // @[Decoder.scala 144:28]
  wire  dram0Handler_io_in_ready; // @[Decoder.scala 144:28]
  wire  dram0Handler_io_in_valid; // @[Decoder.scala 144:28]
  wire  dram0Handler_io_in_bits_write; // @[Decoder.scala 144:28]
  wire [20:0] dram0Handler_io_in_bits_address; // @[Decoder.scala 144:28]
  wire [20:0] dram0Handler_io_in_bits_size; // @[Decoder.scala 144:28]
  wire [2:0] dram0Handler_io_in_bits_stride; // @[Decoder.scala 144:28]
  wire  dram0Handler_io_in_bits_reverse; // @[Decoder.scala 144:28]
  wire  dram0Handler_io_out_ready; // @[Decoder.scala 144:28]
  wire  dram0Handler_io_out_valid; // @[Decoder.scala 144:28]
  wire  dram0Handler_io_out_bits_write; // @[Decoder.scala 144:28]
  wire [20:0] dram0Handler_io_out_bits_address; // @[Decoder.scala 144:28]
  wire [20:0] dram0Handler_io_out_bits_size; // @[Decoder.scala 144:28]
  wire  dram1Handler_clock; // @[Decoder.scala 153:28]
  wire  dram1Handler_reset; // @[Decoder.scala 153:28]
  wire  dram1Handler_io_in_ready; // @[Decoder.scala 153:28]
  wire  dram1Handler_io_in_valid; // @[Decoder.scala 153:28]
  wire  dram1Handler_io_in_bits_write; // @[Decoder.scala 153:28]
  wire [20:0] dram1Handler_io_in_bits_address; // @[Decoder.scala 153:28]
  wire [20:0] dram1Handler_io_in_bits_size; // @[Decoder.scala 153:28]
  wire [2:0] dram1Handler_io_in_bits_stride; // @[Decoder.scala 153:28]
  wire  dram1Handler_io_in_bits_reverse; // @[Decoder.scala 153:28]
  wire  dram1Handler_io_out_ready; // @[Decoder.scala 153:28]
  wire  dram1Handler_io_out_valid; // @[Decoder.scala 153:28]
  wire  dram1Handler_io_out_bits_write; // @[Decoder.scala 153:28]
  wire [20:0] dram1Handler_io_out_bits_address; // @[Decoder.scala 153:28]
  wire [20:0] dram1Handler_io_out_bits_size; // @[Decoder.scala 153:28]
  wire  dram0_clock; // @[Mem.scala 22:19]
  wire  dram0_reset; // @[Mem.scala 22:19]
  wire  dram0_io_enq_ready; // @[Mem.scala 22:19]
  wire  dram0_io_enq_valid; // @[Mem.scala 22:19]
  wire  dram0_io_enq_bits_write; // @[Mem.scala 22:19]
  wire [20:0] dram0_io_enq_bits_address; // @[Mem.scala 22:19]
  wire [20:0] dram0_io_enq_bits_size; // @[Mem.scala 22:19]
  wire [2:0] dram0_io_enq_bits_stride; // @[Mem.scala 22:19]
  wire  dram0_io_deq_ready; // @[Mem.scala 22:19]
  wire  dram0_io_deq_valid; // @[Mem.scala 22:19]
  wire  dram0_io_deq_bits_write; // @[Mem.scala 22:19]
  wire [20:0] dram0_io_deq_bits_address; // @[Mem.scala 22:19]
  wire [20:0] dram0_io_deq_bits_size; // @[Mem.scala 22:19]
  wire [2:0] dram0_io_deq_bits_stride; // @[Mem.scala 22:19]
  wire  dram0_io_deq_bits_reverse; // @[Mem.scala 22:19]
  wire  dram1_clock; // @[Mem.scala 22:19]
  wire  dram1_reset; // @[Mem.scala 22:19]
  wire  dram1_io_enq_ready; // @[Mem.scala 22:19]
  wire  dram1_io_enq_valid; // @[Mem.scala 22:19]
  wire  dram1_io_enq_bits_write; // @[Mem.scala 22:19]
  wire [20:0] dram1_io_enq_bits_address; // @[Mem.scala 22:19]
  wire [20:0] dram1_io_enq_bits_size; // @[Mem.scala 22:19]
  wire [2:0] dram1_io_enq_bits_stride; // @[Mem.scala 22:19]
  wire  dram1_io_deq_ready; // @[Mem.scala 22:19]
  wire  dram1_io_deq_valid; // @[Mem.scala 22:19]
  wire  dram1_io_deq_bits_write; // @[Mem.scala 22:19]
  wire [20:0] dram1_io_deq_bits_address; // @[Mem.scala 22:19]
  wire [20:0] dram1_io_deq_bits_size; // @[Mem.scala 22:19]
  wire [2:0] dram1_io_deq_bits_stride; // @[Mem.scala 22:19]
  wire  dram1_io_deq_bits_reverse; // @[Mem.scala 22:19]
  wire  memPortAHandler_clock; // @[Decoder.scala 168:31]
  wire  memPortAHandler_reset; // @[Decoder.scala 168:31]
  wire  memPortAHandler_io_in_ready; // @[Decoder.scala 168:31]
  wire  memPortAHandler_io_in_valid; // @[Decoder.scala 168:31]
  wire  memPortAHandler_io_in_bits_write; // @[Decoder.scala 168:31]
  wire [13:0] memPortAHandler_io_in_bits_address; // @[Decoder.scala 168:31]
  wire [13:0] memPortAHandler_io_in_bits_size; // @[Decoder.scala 168:31]
  wire [2:0] memPortAHandler_io_in_bits_stride; // @[Decoder.scala 168:31]
  wire  memPortAHandler_io_in_bits_reverse; // @[Decoder.scala 168:31]
  wire  memPortAHandler_io_out_ready; // @[Decoder.scala 168:31]
  wire  memPortAHandler_io_out_valid; // @[Decoder.scala 168:31]
  wire  memPortAHandler_io_out_bits_write; // @[Decoder.scala 168:31]
  wire [13:0] memPortAHandler_io_out_bits_address; // @[Decoder.scala 168:31]
  wire  memPortBHandler_clock; // @[Decoder.scala 177:31]
  wire  memPortBHandler_reset; // @[Decoder.scala 177:31]
  wire  memPortBHandler_io_in_ready; // @[Decoder.scala 177:31]
  wire  memPortBHandler_io_in_valid; // @[Decoder.scala 177:31]
  wire  memPortBHandler_io_in_bits_write; // @[Decoder.scala 177:31]
  wire [13:0] memPortBHandler_io_in_bits_address; // @[Decoder.scala 177:31]
  wire [13:0] memPortBHandler_io_in_bits_size; // @[Decoder.scala 177:31]
  wire [2:0] memPortBHandler_io_in_bits_stride; // @[Decoder.scala 177:31]
  wire  memPortBHandler_io_in_bits_reverse; // @[Decoder.scala 177:31]
  wire  memPortBHandler_io_out_ready; // @[Decoder.scala 177:31]
  wire  memPortBHandler_io_out_valid; // @[Decoder.scala 177:31]
  wire  memPortBHandler_io_out_bits_write; // @[Decoder.scala 177:31]
  wire [13:0] memPortBHandler_io_out_bits_address; // @[Decoder.scala 177:31]
  wire  lockPool_clock; // @[Decoder.scala 193:24]
  wire  lockPool_reset; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_0_in_ready; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_0_in_valid; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_0_in_bits_write; // @[Decoder.scala 193:24]
  wire [13:0] lockPool_io_actor_0_in_bits_address; // @[Decoder.scala 193:24]
  wire [13:0] lockPool_io_actor_0_in_bits_size; // @[Decoder.scala 193:24]
  wire [2:0] lockPool_io_actor_0_in_bits_stride; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_0_in_bits_reverse; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_0_out_ready; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_0_out_valid; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_0_out_bits_write; // @[Decoder.scala 193:24]
  wire [13:0] lockPool_io_actor_0_out_bits_address; // @[Decoder.scala 193:24]
  wire [13:0] lockPool_io_actor_0_out_bits_size; // @[Decoder.scala 193:24]
  wire [2:0] lockPool_io_actor_0_out_bits_stride; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_0_out_bits_reverse; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_1_in_ready; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_1_in_valid; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_1_in_bits_write; // @[Decoder.scala 193:24]
  wire [13:0] lockPool_io_actor_1_in_bits_address; // @[Decoder.scala 193:24]
  wire [13:0] lockPool_io_actor_1_in_bits_size; // @[Decoder.scala 193:24]
  wire [2:0] lockPool_io_actor_1_in_bits_stride; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_1_out_ready; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_1_out_valid; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_1_out_bits_write; // @[Decoder.scala 193:24]
  wire [13:0] lockPool_io_actor_1_out_bits_address; // @[Decoder.scala 193:24]
  wire [13:0] lockPool_io_actor_1_out_bits_size; // @[Decoder.scala 193:24]
  wire [2:0] lockPool_io_actor_1_out_bits_stride; // @[Decoder.scala 193:24]
  wire  lockPool_io_actor_1_out_bits_reverse; // @[Decoder.scala 193:24]
  wire  lockPool_io_lock_ready; // @[Decoder.scala 193:24]
  wire  lockPool_io_lock_valid; // @[Decoder.scala 193:24]
  wire  lockPool_io_lock_bits_cond_write; // @[Decoder.scala 193:24]
  wire [13:0] lockPool_io_lock_bits_cond_address; // @[Decoder.scala 193:24]
  wire [13:0] lockPool_io_lock_bits_cond_size; // @[Decoder.scala 193:24]
  wire [2:0] lockPool_io_lock_bits_cond_stride; // @[Decoder.scala 193:24]
  wire  lockPool_io_lock_bits_cond_reverse; // @[Decoder.scala 193:24]
  wire  lockPool_io_lock_bits_lock; // @[Decoder.scala 193:24]
  wire  lockPool_io_lock_bits_by; // @[Decoder.scala 193:24]
  wire  accHandler_clock; // @[Decoder.scala 207:26]
  wire  accHandler_reset; // @[Decoder.scala 207:26]
  wire  accHandler_io_in_ready; // @[Decoder.scala 207:26]
  wire  accHandler_io_in_valid; // @[Decoder.scala 207:26]
  wire [3:0] accHandler_io_in_bits_instruction_op; // @[Decoder.scala 207:26]
  wire  accHandler_io_in_bits_instruction_sourceLeft; // @[Decoder.scala 207:26]
  wire  accHandler_io_in_bits_instruction_sourceRight; // @[Decoder.scala 207:26]
  wire  accHandler_io_in_bits_instruction_dest; // @[Decoder.scala 207:26]
  wire [11:0] accHandler_io_in_bits_address; // @[Decoder.scala 207:26]
  wire [11:0] accHandler_io_in_bits_altAddress; // @[Decoder.scala 207:26]
  wire  accHandler_io_in_bits_read; // @[Decoder.scala 207:26]
  wire  accHandler_io_in_bits_write; // @[Decoder.scala 207:26]
  wire  accHandler_io_in_bits_accumulate; // @[Decoder.scala 207:26]
  wire [11:0] accHandler_io_in_bits_size; // @[Decoder.scala 207:26]
  wire [2:0] accHandler_io_in_bits_stride; // @[Decoder.scala 207:26]
  wire  accHandler_io_in_bits_reverse; // @[Decoder.scala 207:26]
  wire  accHandler_io_out_ready; // @[Decoder.scala 207:26]
  wire  accHandler_io_out_valid; // @[Decoder.scala 207:26]
  wire [3:0] accHandler_io_out_bits_instruction_op; // @[Decoder.scala 207:26]
  wire  accHandler_io_out_bits_instruction_sourceLeft; // @[Decoder.scala 207:26]
  wire  accHandler_io_out_bits_instruction_sourceRight; // @[Decoder.scala 207:26]
  wire  accHandler_io_out_bits_instruction_dest; // @[Decoder.scala 207:26]
  wire [11:0] accHandler_io_out_bits_address; // @[Decoder.scala 207:26]
  wire [11:0] accHandler_io_out_bits_altAddress; // @[Decoder.scala 207:26]
  wire  accHandler_io_out_bits_read; // @[Decoder.scala 207:26]
  wire  accHandler_io_out_bits_write; // @[Decoder.scala 207:26]
  wire  accHandler_io_out_bits_accumulate; // @[Decoder.scala 207:26]
  wire  acc_clock; // @[Mem.scala 22:19]
  wire  acc_reset; // @[Mem.scala 22:19]
  wire  acc_io_enq_ready; // @[Mem.scala 22:19]
  wire  acc_io_enq_valid; // @[Mem.scala 22:19]
  wire [3:0] acc_io_enq_bits_instruction_op; // @[Mem.scala 22:19]
  wire  acc_io_enq_bits_instruction_sourceLeft; // @[Mem.scala 22:19]
  wire  acc_io_enq_bits_instruction_sourceRight; // @[Mem.scala 22:19]
  wire  acc_io_enq_bits_instruction_dest; // @[Mem.scala 22:19]
  wire [11:0] acc_io_enq_bits_address; // @[Mem.scala 22:19]
  wire [11:0] acc_io_enq_bits_altAddress; // @[Mem.scala 22:19]
  wire  acc_io_enq_bits_read; // @[Mem.scala 22:19]
  wire  acc_io_enq_bits_write; // @[Mem.scala 22:19]
  wire  acc_io_enq_bits_accumulate; // @[Mem.scala 22:19]
  wire [11:0] acc_io_enq_bits_size; // @[Mem.scala 22:19]
  wire [2:0] acc_io_enq_bits_stride; // @[Mem.scala 22:19]
  wire  acc_io_deq_ready; // @[Mem.scala 22:19]
  wire  acc_io_deq_valid; // @[Mem.scala 22:19]
  wire [3:0] acc_io_deq_bits_instruction_op; // @[Mem.scala 22:19]
  wire  acc_io_deq_bits_instruction_sourceLeft; // @[Mem.scala 22:19]
  wire  acc_io_deq_bits_instruction_sourceRight; // @[Mem.scala 22:19]
  wire  acc_io_deq_bits_instruction_dest; // @[Mem.scala 22:19]
  wire [11:0] acc_io_deq_bits_address; // @[Mem.scala 22:19]
  wire [11:0] acc_io_deq_bits_altAddress; // @[Mem.scala 22:19]
  wire  acc_io_deq_bits_read; // @[Mem.scala 22:19]
  wire  acc_io_deq_bits_write; // @[Mem.scala 22:19]
  wire  acc_io_deq_bits_accumulate; // @[Mem.scala 22:19]
  wire [11:0] acc_io_deq_bits_size; // @[Mem.scala 22:19]
  wire [2:0] acc_io_deq_bits_stride; // @[Mem.scala 22:19]
  wire  acc_io_deq_bits_reverse; // @[Mem.scala 22:19]
  wire  arrayHandler_clock; // @[Decoder.scala 230:28]
  wire  arrayHandler_reset; // @[Decoder.scala 230:28]
  wire  arrayHandler_io_in_ready; // @[Decoder.scala 230:28]
  wire  arrayHandler_io_in_valid; // @[Decoder.scala 230:28]
  wire  arrayHandler_io_in_bits_load; // @[Decoder.scala 230:28]
  wire  arrayHandler_io_in_bits_zeroes; // @[Decoder.scala 230:28]
  wire [13:0] arrayHandler_io_in_bits_size; // @[Decoder.scala 230:28]
  wire  arrayHandler_io_out_ready; // @[Decoder.scala 230:28]
  wire  arrayHandler_io_out_valid; // @[Decoder.scala 230:28]
  wire  arrayHandler_io_out_bits_load; // @[Decoder.scala 230:28]
  wire  arrayHandler_io_out_bits_zeroes; // @[Decoder.scala 230:28]
  wire  array_clock; // @[Mem.scala 22:19]
  wire  array_reset; // @[Mem.scala 22:19]
  wire  array_io_enq_ready; // @[Mem.scala 22:19]
  wire  array_io_enq_valid; // @[Mem.scala 22:19]
  wire  array_io_enq_bits_load; // @[Mem.scala 22:19]
  wire  array_io_enq_bits_zeroes; // @[Mem.scala 22:19]
  wire [13:0] array_io_enq_bits_size; // @[Mem.scala 22:19]
  wire  array_io_deq_ready; // @[Mem.scala 22:19]
  wire  array_io_deq_valid; // @[Mem.scala 22:19]
  wire  array_io_deq_bits_load; // @[Mem.scala 22:19]
  wire  array_io_deq_bits_zeroes; // @[Mem.scala 22:19]
  wire [13:0] array_io_deq_bits_size; // @[Mem.scala 22:19]
  wire  dataflow_clock; // @[Mem.scala 22:19]
  wire  dataflow_reset; // @[Mem.scala 22:19]
  wire  dataflow_io_enq_ready; // @[Mem.scala 22:19]
  wire  dataflow_io_enq_valid; // @[Mem.scala 22:19]
  wire [3:0] dataflow_io_enq_bits_kind; // @[Mem.scala 22:19]
  wire [13:0] dataflow_io_enq_bits_size; // @[Mem.scala 22:19]
  wire  dataflow_io_deq_ready; // @[Mem.scala 22:19]
  wire  dataflow_io_deq_valid; // @[Mem.scala 22:19]
  wire [3:0] dataflow_io_deq_bits_kind; // @[Mem.scala 22:19]
  wire [13:0] dataflow_io_deq_bits_size; // @[Mem.scala 22:19]
  wire  hostDataflowHandler_clock; // @[Decoder.scala 250:35]
  wire  hostDataflowHandler_reset; // @[Decoder.scala 250:35]
  wire  hostDataflowHandler_io_in_ready; // @[Decoder.scala 250:35]
  wire  hostDataflowHandler_io_in_valid; // @[Decoder.scala 250:35]
  wire [1:0] hostDataflowHandler_io_in_bits_kind; // @[Decoder.scala 250:35]
  wire [13:0] hostDataflowHandler_io_in_bits_size; // @[Decoder.scala 250:35]
  wire  hostDataflowHandler_io_out_ready; // @[Decoder.scala 250:35]
  wire  hostDataflowHandler_io_out_valid; // @[Decoder.scala 250:35]
  wire [1:0] hostDataflowHandler_io_out_bits_kind; // @[Decoder.scala 250:35]
  wire  hostDataflow_clock; // @[Mem.scala 22:19]
  wire  hostDataflow_reset; // @[Mem.scala 22:19]
  wire  hostDataflow_io_enq_ready; // @[Mem.scala 22:19]
  wire  hostDataflow_io_enq_valid; // @[Mem.scala 22:19]
  wire [1:0] hostDataflow_io_enq_bits_kind; // @[Mem.scala 22:19]
  wire [13:0] hostDataflow_io_enq_bits_size; // @[Mem.scala 22:19]
  wire  hostDataflow_io_deq_ready; // @[Mem.scala 22:19]
  wire  hostDataflow_io_deq_valid; // @[Mem.scala 22:19]
  wire [1:0] hostDataflow_io_deq_bits_kind; // @[Mem.scala 22:19]
  wire [13:0] hostDataflow_io_deq_bits_size; // @[Mem.scala 22:19]
  wire  enqueuer1_clock; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer1_reset; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer1_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer1_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer1_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer1_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_clock; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_reset; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer3_clock; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer3_reset; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer3_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer3_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer3_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer3_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer3_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer3_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer3_io_out_2_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer3_io_out_2_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_clock; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_reset; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_io_out_2_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_io_out_2_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_io_out_3_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer4_io_out_3_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_clock; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_reset; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_out_2_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_out_2_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_out_3_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_out_3_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_out_4_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer5_io_out_4_valid; // @[MultiEnqueue.scala 182:43]
  reg [15:0] timeout; // @[Decoder.scala 96:24]
  reg [15:0] timer; // @[Decoder.scala 97:24]
  wire [15:0] _timer_T_1 = timer + 16'h1; // @[Decoder.scala 102:22]
  reg [31:0] tracepoint; // @[Decoder.scala 108:31]
  reg [31:0] programCounter; // @[Decoder.scala 109:31]
  wire [31:0] _programCounter_T_1 = programCounter + 32'h1; // @[Decoder.scala 111:38]
  wire [31:0] _GEN_2 = instruction_io_deq_ready & instruction_io_deq_valid ? _programCounter_T_1 : programCounter; // @[Decoder.scala 110:48 111:20 109:31]
  reg [31:0] dram0AddressOffset; // @[Decoder.scala 126:35]
  reg [3:0] dram0CacheBehaviour; // @[Decoder.scala 129:36]
  reg [31:0] dram1AddressOffset; // @[Decoder.scala 130:35]
  reg [3:0] dram1CacheBehaviour; // @[Decoder.scala 133:36]
  wire  io_acc_bits_isMemControl = accHandler_io_out_bits_instruction_op == 4'h0; // @[AccumulatorWithALUArrayControl.scala 101:39]
  wire [11:0] _GEN_3 = accHandler_io_out_bits_write ? accHandler_io_out_bits_altAddress : accHandler_io_out_bits_address
    ; // @[AccumulatorWithALUArrayControl.scala 111:21 112:25 115:25]
  wire [11:0] _GEN_4 = accHandler_io_out_bits_write ? accHandler_io_out_bits_address : accHandler_io_out_bits_altAddress
    ; // @[AccumulatorWithALUArrayControl.scala 111:21 113:26 116:26]
  wire [11:0] _GEN_5 = accHandler_io_out_bits_read ? accHandler_io_out_bits_address : _GEN_3; // @[AccumulatorWithALUArrayControl.scala 107:18 108:23]
  wire [11:0] _GEN_6 = accHandler_io_out_bits_read ? accHandler_io_out_bits_altAddress : _GEN_4; // @[AccumulatorWithALUArrayControl.scala 107:18 109:24]
  wire [3:0] _flags_WIRE_1 = instruction_io_deq_bits_flags;
  wire  flags_accumulate = _flags_WIRE_1[0]; // @[Decoder.scala 288:45]
  wire  flags_zeroes = _flags_WIRE_1[1]; // @[Decoder.scala 288:45]
  wire [63:0] _args_WIRE_1 = instruction_io_deq_bits_arguments;
  wire [13:0] args_memAddress = _args_WIRE_1[13:0]; // @[Decoder.scala 289:48]
  wire [2:0] args_memStride = _args_WIRE_1[16:14]; // @[Decoder.scala 289:48]
  wire [20:0] args_accAddress = _args_WIRE_1[44:24]; // @[Decoder.scala 289:48]
  wire [2:0] args_accStride = _args_WIRE_1[47:45]; // @[Decoder.scala 289:48]
  wire [15:0] args_size = _args_WIRE_1[63:48]; // @[Decoder.scala 289:48]
  wire [13:0] _instruction_io_deq_ready_w_lock_T = args_memAddress / 14'h2000; // @[Decoder.scala 191:15]
  wire  _GEN_9 = flags_zeroes & instruction_io_deq_valid; // @[Decoder.scala 291:24 MultiEnqueue.scala 114:17 40:17]
  wire  instruction_io_deq_ready_dataflow_io_enq_w_ready = dataflow_io_enq_ready; // @[MultiEnqueue.scala 115:10 ReadyValid.scala 16:17]
  wire  _GEN_10 = flags_zeroes & instruction_io_deq_ready_dataflow_io_enq_w_ready; // @[Decoder.scala 291:24 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  instruction_io_deq_ready_dataflow_io_enq_w_valid = enqueuer3_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  instruction_io_deq_ready_dataflow_io_enq_w_1_valid = enqueuer5_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_11 = flags_zeroes ? instruction_io_deq_ready_dataflow_io_enq_w_valid :
    instruction_io_deq_ready_dataflow_io_enq_w_1_valid; // @[Decoder.scala 291:24 MultiEnqueue.scala 115:10 172:10]
  wire [3:0] _GEN_12 = flags_zeroes ? 4'h3 : 4'h2; // @[Decoder.scala 291:24 MultiEnqueue.scala 115:10 172:10]
  wire [13:0] instruction_io_deq_ready_w_size = args_size[13:0]; // @[Decoder.scala 733:17 735:12]
  wire [13:0] _GEN_13 = flags_zeroes ? instruction_io_deq_ready_w_size : instruction_io_deq_ready_w_size; // @[Decoder.scala 291:24 MultiEnqueue.scala 115:10 172:10]
  wire  instruction_io_deq_ready_array_io_enq_w_ready = array_io_enq_ready; // @[MultiEnqueue.scala 116:10 ReadyValid.scala 16:17]
  wire  _GEN_14 = flags_zeroes & instruction_io_deq_ready_array_io_enq_w_ready; // @[Decoder.scala 291:24 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  instruction_io_deq_ready_array_io_enq_w_valid = enqueuer3_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  instruction_io_deq_ready_array_io_enq_w_1_valid = enqueuer5_io_out_2_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_15 = flags_zeroes ? instruction_io_deq_ready_array_io_enq_w_valid :
    instruction_io_deq_ready_array_io_enq_w_1_valid; // @[Decoder.scala 291:24 MultiEnqueue.scala 116:10 174:10]
  wire  instruction_io_deq_ready_acc_io_enq_w_ready = acc_io_enq_ready; // @[MultiEnqueue.scala 117:10 ReadyValid.scala 16:17]
  wire  _GEN_19 = flags_zeroes & instruction_io_deq_ready_acc_io_enq_w_ready; // @[Decoder.scala 291:24 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  instruction_io_deq_ready_acc_io_enq_w_valid = enqueuer3_io_out_2_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  instruction_io_deq_ready_acc_io_enq_w_1_valid = enqueuer5_io_out_3_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_20 = flags_zeroes ? instruction_io_deq_ready_acc_io_enq_w_valid :
    instruction_io_deq_ready_acc_io_enq_w_1_valid; // @[Decoder.scala 291:24 MultiEnqueue.scala 117:10 175:10]
  wire [11:0] instruction_io_deq_ready_w_2_address = args_accAddress[11:0]; // @[Decoder.scala 716:17 718:15]
  wire [11:0] _GEN_25 = flags_zeroes ? instruction_io_deq_ready_w_2_address : instruction_io_deq_ready_w_2_address; // @[Decoder.scala 291:24 MultiEnqueue.scala 117:10 175:10]
  wire [11:0] instruction_io_deq_ready_w_2_size = args_size[11:0]; // @[Decoder.scala 716:17 723:12]
  wire [11:0] _GEN_30 = flags_zeroes ? instruction_io_deq_ready_w_2_size : instruction_io_deq_ready_w_2_size; // @[Decoder.scala 291:24 MultiEnqueue.scala 117:10 175:10]
  wire  _GEN_33 = flags_zeroes ? enqueuer3_io_in_ready : enqueuer5_io_in_ready; // @[Decoder.scala 291:24 292:25 314:25]
  wire  _GEN_34 = flags_zeroes ? 1'h0 : instruction_io_deq_valid; // @[Decoder.scala 291:24 MultiEnqueue.scala 171:17 40:17]
  wire  _GEN_35 = flags_zeroes ? 1'h0 : instruction_io_deq_ready_dataflow_io_enq_w_ready; // @[Decoder.scala 291:24 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  instruction_io_deq_ready_lockPool_io_actor_0_in_w_ready = lockPool_io_actor_0_in_ready; // @[ReadyValid.scala 16:17 MultiEnqueue.scala 173:10]
  wire  _GEN_36 = flags_zeroes ? 1'h0 : instruction_io_deq_ready_lockPool_io_actor_0_in_w_ready; // @[Decoder.scala 291:24 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  instruction_io_deq_ready_lockPool_io_actor_0_in_w_valid = enqueuer5_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_37 = flags_zeroes ? 1'h0 : instruction_io_deq_ready_lockPool_io_actor_0_in_w_valid; // @[Decoder.scala 291:24 670:16 MultiEnqueue.scala 173:10]
  wire [13:0] _GEN_39 = flags_zeroes ? 14'h0 : args_memAddress; // @[Decoder.scala 291:24 669:15 MultiEnqueue.scala 173:10]
  wire [13:0] _GEN_40 = flags_zeroes ? 14'h0 : instruction_io_deq_ready_w_size; // @[Decoder.scala 291:24 669:15 MultiEnqueue.scala 173:10]
  wire [2:0] _GEN_41 = flags_zeroes ? 3'h0 : args_memStride; // @[Decoder.scala 291:24 669:15 MultiEnqueue.scala 173:10]
  wire  _GEN_43 = flags_zeroes ? 1'h0 : instruction_io_deq_ready_array_io_enq_w_ready; // @[Decoder.scala 291:24 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  _GEN_44 = flags_zeroes ? 1'h0 : instruction_io_deq_ready_acc_io_enq_w_ready; // @[Decoder.scala 291:24 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  instruction_io_deq_ready_lockPool_io_lock_w_ready = lockPool_io_lock_ready; // @[ReadyValid.scala 16:17 MultiEnqueue.scala 176:10]
  wire  _GEN_45 = flags_zeroes ? 1'h0 : instruction_io_deq_ready_lockPool_io_lock_w_ready; // @[Decoder.scala 291:24 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  instruction_io_deq_ready_lockPool_io_lock_w_valid = enqueuer5_io_out_4_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_46 = flags_zeroes ? 1'h0 : instruction_io_deq_ready_lockPool_io_lock_w_valid; // @[Decoder.scala 291:24 Decoupled.scala 72:20 MultiEnqueue.scala 176:10]
  wire  instruction_io_deq_ready_w_6_lock = _instruction_io_deq_ready_w_lock_T[0]; // @[Decoder.scala 755:17 758:12]
  wire  _T_3 = instruction_io_deq_bits_opcode == 4'h3; // @[Decoder.scala 333:38]
  wire [13:0] args_1_address = instruction_io_deq_bits_arguments[13:0]; // @[Decoder.scala 341:48]
  wire [2:0] args_1_stride = instruction_io_deq_bits_arguments[16:14]; // @[Decoder.scala 341:48]
  wire [23:0] args_1_size = instruction_io_deq_bits_arguments[47:24]; // @[Decoder.scala 341:48]
  wire [7:0] stride = 8'h1 << args_1_stride; // @[Decoder.scala 350:24]
  wire [31:0] _req_T = args_1_size * stride; // @[Decoder.scala 352:35]
  wire [31:0] _GEN_55 = {{18'd0}, args_1_address}; // @[Decoder.scala 352:22]
  wire [31:0] _req_T_2 = _GEN_55 + _req_T; // @[Decoder.scala 352:22]
  wire [13:0] req_1_address = _req_T_2[13:0]; // @[MemControl.scala 44:19 45:17]
  wire [13:0] _instruction_io_deq_ready_w_lock_T_1 = req_1_address / 14'h2000; // @[Decoder.scala 191:15]
  wire  _GEN_56 = flags_accumulate & instruction_io_deq_valid; // @[Decoder.scala 343:24 MultiEnqueue.scala 40:17 60:17]
  wire  _GEN_57 = flags_accumulate & instruction_io_deq_ready_array_io_enq_w_ready; // @[Decoder.scala 343:24 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  instruction_io_deq_ready_array_io_enq_w_2_valid = enqueuer1_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  instruction_io_deq_ready_array_io_enq_w_3_valid = enqueuer4_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_58 = flags_accumulate ? instruction_io_deq_ready_array_io_enq_w_2_valid :
    instruction_io_deq_ready_array_io_enq_w_3_valid; // @[Decoder.scala 343:24 MultiEnqueue.scala 152:10 61:10]
  wire [13:0] instruction_io_deq_ready_w_7_size = args_1_size[13:0]; // @[Decoder.scala 744:17 747:12]
  wire [13:0] _GEN_61 = flags_accumulate ? instruction_io_deq_ready_w_7_size : instruction_io_deq_ready_w_7_size; // @[Decoder.scala 343:24 MultiEnqueue.scala 152:10 61:10]
  wire  _GEN_62 = flags_accumulate ? enqueuer1_io_in_ready : enqueuer4_io_in_ready; // @[Decoder.scala 343:24 344:25 358:25]
  wire  _GEN_63 = flags_accumulate ? 1'h0 : instruction_io_deq_valid; // @[Decoder.scala 343:24 MultiEnqueue.scala 150:17 40:17]
  wire  _GEN_64 = flags_accumulate ? 1'h0 : instruction_io_deq_ready_dataflow_io_enq_w_ready; // @[Decoder.scala 343:24 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  instruction_io_deq_ready_dataflow_io_enq_w_2_valid = enqueuer4_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_65 = flags_accumulate ? 1'h0 : instruction_io_deq_ready_dataflow_io_enq_w_2_valid; // @[Decoder.scala 343:24 670:16 MultiEnqueue.scala 151:10]
  wire [3:0] _GEN_66 = flags_accumulate ? 4'h0 : 4'h1; // @[Decoder.scala 343:24 669:15 MultiEnqueue.scala 151:10]
  wire [13:0] _GEN_67 = flags_accumulate ? 14'h0 : instruction_io_deq_ready_w_7_size; // @[Decoder.scala 343:24 669:15 MultiEnqueue.scala 151:10]
  wire  _GEN_68 = flags_accumulate ? 1'h0 : instruction_io_deq_ready_array_io_enq_w_ready; // @[Decoder.scala 343:24 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  _GEN_69 = flags_accumulate ? 1'h0 : instruction_io_deq_ready_lockPool_io_actor_0_in_w_ready; // @[Decoder.scala 343:24 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  instruction_io_deq_ready_lockPool_io_actor_0_in_w_1_valid = enqueuer4_io_out_2_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_70 = flags_accumulate ? 1'h0 : instruction_io_deq_ready_lockPool_io_actor_0_in_w_1_valid; // @[Decoder.scala 343:24 670:16 MultiEnqueue.scala 153:10]
  wire [13:0] _GEN_72 = flags_accumulate ? 14'h0 : req_1_address; // @[Decoder.scala 343:24 669:15 MultiEnqueue.scala 153:10]
  wire [2:0] _GEN_74 = flags_accumulate ? 3'h0 : args_1_stride; // @[Decoder.scala 343:24 669:15 MultiEnqueue.scala 153:10]
  wire  _GEN_75 = flags_accumulate ? 1'h0 : 1'h1; // @[Decoder.scala 343:24 669:15 MultiEnqueue.scala 153:10]
  wire  _GEN_76 = flags_accumulate ? 1'h0 : instruction_io_deq_ready_lockPool_io_lock_w_ready; // @[Decoder.scala 343:24 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  instruction_io_deq_ready_lockPool_io_lock_w_1_valid = enqueuer4_io_out_3_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_77 = flags_accumulate ? 1'h0 : instruction_io_deq_ready_lockPool_io_lock_w_1_valid; // @[Decoder.scala 343:24 Decoupled.scala 72:20 MultiEnqueue.scala 154:10]
  wire  instruction_io_deq_ready_w_10_lock = _instruction_io_deq_ready_w_lock_T_1[0]; // @[Decoder.scala 755:17 758:12]
  wire  _T_6 = _flags_WIRE_1 == 4'h1; // @[Decoder.scala 412:27]
  wire  _T_7 = _flags_WIRE_1 == 4'h2; // @[Decoder.scala 441:27]
  wire  _T_8 = _flags_WIRE_1 == 4'h3; // @[Decoder.scala 470:27]
  wire  _T_9 = _flags_WIRE_1 == 4'hc; // @[Decoder.scala 499:18]
  wire  _T_10 = _flags_WIRE_1 == 4'hd; // @[Decoder.scala 524:18]
  wire  _T_11 = _flags_WIRE_1 == 4'hf; // @[Decoder.scala 549:18]
  wire  _GEN_87 = _T_11 & instruction_io_deq_valid; // @[Decoder.scala 550:7 MultiEnqueue.scala 150:17 40:17]
  wire  _GEN_88 = _T_11 & instruction_io_deq_ready_dataflow_io_enq_w_ready; // @[Decoder.scala 550:7 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  _GEN_89 = _T_11 & instruction_io_deq_ready_dataflow_io_enq_w_2_valid; // @[Decoder.scala 550:7 MultiEnqueue.scala 151:10 Decoder.scala 670:16]
  wire [3:0] _GEN_90 = _T_11 ? 4'h5 : 4'h0; // @[Decoder.scala 550:7 MultiEnqueue.scala 151:10 Decoder.scala 669:15]
  wire [13:0] _GEN_91 = _T_11 ? instruction_io_deq_ready_w_size : 14'h0; // @[Decoder.scala 550:7 MultiEnqueue.scala 151:10 Decoder.scala 669:15]
  wire  _GEN_92 = _T_11 & instruction_io_deq_ready_lockPool_io_actor_0_in_w_ready; // @[Decoder.scala 550:7 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  _GEN_93 = _T_11 & instruction_io_deq_ready_array_io_enq_w_3_valid; // @[Decoder.scala 550:7 MultiEnqueue.scala 152:10 Decoder.scala 670:16]
  wire [13:0] _GEN_95 = _T_11 ? args_memAddress : 14'h0; // @[Decoder.scala 550:7 MultiEnqueue.scala 152:10 Decoder.scala 669:15]
  wire [2:0] _GEN_97 = _T_11 ? args_memStride : 3'h0; // @[Decoder.scala 550:7 MultiEnqueue.scala 152:10 Decoder.scala 669:15]
  wire  _GEN_99 = _T_11 & instruction_io_deq_ready_acc_io_enq_w_ready; // @[Decoder.scala 550:7 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  _GEN_100 = _T_11 & instruction_io_deq_ready_lockPool_io_actor_0_in_w_1_valid; // @[Decoder.scala 550:7 MultiEnqueue.scala 153:10 Decoder.scala 670:16]
  wire [11:0] _GEN_105 = _T_11 ? instruction_io_deq_ready_w_2_address : 12'h0; // @[Decoder.scala 550:7 MultiEnqueue.scala 153:10 Decoder.scala 669:15]
  wire [11:0] _GEN_110 = _T_11 ? instruction_io_deq_ready_w_2_size : 12'h0; // @[Decoder.scala 550:7 MultiEnqueue.scala 153:10 Decoder.scala 669:15]
  wire [2:0] _GEN_111 = _T_11 ? args_accStride : 3'h0; // @[Decoder.scala 550:7 MultiEnqueue.scala 153:10 Decoder.scala 669:15]
  wire  _GEN_113 = _T_11 & instruction_io_deq_ready_lockPool_io_lock_w_ready; // @[Decoder.scala 550:7 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  _GEN_114 = _T_11 & instruction_io_deq_ready_lockPool_io_lock_w_1_valid; // @[Decoder.scala 550:7 MultiEnqueue.scala 154:10 Decoupled.scala 72:20]
  wire  _GEN_124 = _T_11 ? enqueuer4_io_in_ready : 1'h1; // @[Decoder.scala 550:7 559:25 575:25]
  wire  _GEN_125 = _T_10 ? instruction_io_deq_valid : _GEN_87; // @[Decoder.scala 525:7 MultiEnqueue.scala 150:17]
  wire  _GEN_126 = _T_10 ? instruction_io_deq_ready_dataflow_io_enq_w_ready : _GEN_88; // @[Decoder.scala 525:7 ReadyValid.scala 19:11]
  wire  _GEN_127 = _T_10 ? instruction_io_deq_ready_dataflow_io_enq_w_2_valid : _GEN_89; // @[Decoder.scala 525:7 MultiEnqueue.scala 151:10]
  wire [3:0] _GEN_128 = _T_10 ? 4'h5 : _GEN_90; // @[Decoder.scala 525:7 MultiEnqueue.scala 151:10]
  wire [13:0] _GEN_129 = _T_10 ? instruction_io_deq_ready_w_size : _GEN_91; // @[Decoder.scala 525:7 MultiEnqueue.scala 151:10]
  wire  _GEN_130 = _T_10 ? instruction_io_deq_ready_lockPool_io_actor_0_in_w_ready : _GEN_92; // @[Decoder.scala 525:7 ReadyValid.scala 19:11]
  wire  _GEN_131 = _T_10 ? instruction_io_deq_ready_array_io_enq_w_3_valid : _GEN_93; // @[Decoder.scala 525:7 MultiEnqueue.scala 152:10]
  wire [13:0] _GEN_133 = _T_10 ? args_memAddress : _GEN_95; // @[Decoder.scala 525:7 MultiEnqueue.scala 152:10]
  wire [2:0] _GEN_135 = _T_10 ? args_memStride : _GEN_97; // @[Decoder.scala 525:7 MultiEnqueue.scala 152:10]
  wire  _GEN_137 = _T_10 ? instruction_io_deq_ready_acc_io_enq_w_ready : _GEN_99; // @[Decoder.scala 525:7 ReadyValid.scala 19:11]
  wire  _GEN_138 = _T_10 ? instruction_io_deq_ready_lockPool_io_actor_0_in_w_1_valid : _GEN_100; // @[Decoder.scala 525:7 MultiEnqueue.scala 153:10]
  wire [11:0] _GEN_143 = _T_10 ? instruction_io_deq_ready_w_2_address : _GEN_105; // @[Decoder.scala 525:7 MultiEnqueue.scala 153:10]
  wire  _GEN_146 = _T_10 | _T_11; // @[Decoder.scala 525:7 MultiEnqueue.scala 153:10]
  wire  _GEN_147 = _T_10 ? 1'h0 : _T_11; // @[Decoder.scala 525:7 MultiEnqueue.scala 153:10]
  wire [11:0] _GEN_148 = _T_10 ? instruction_io_deq_ready_w_2_size : _GEN_110; // @[Decoder.scala 525:7 MultiEnqueue.scala 153:10]
  wire [2:0] _GEN_149 = _T_10 ? args_accStride : _GEN_111; // @[Decoder.scala 525:7 MultiEnqueue.scala 153:10]
  wire  _GEN_151 = _T_10 ? instruction_io_deq_ready_lockPool_io_lock_w_ready : _GEN_113; // @[Decoder.scala 525:7 ReadyValid.scala 19:11]
  wire  _GEN_152 = _T_10 ? instruction_io_deq_ready_lockPool_io_lock_w_1_valid : _GEN_114; // @[Decoder.scala 525:7 MultiEnqueue.scala 154:10]
  wire [13:0] _GEN_155 = _T_10 ? instruction_io_deq_ready_w_size : instruction_io_deq_ready_w_size; // @[Decoder.scala 525:7 MultiEnqueue.scala 154:10]
  wire  _GEN_158 = _T_10 ? instruction_io_deq_ready_w_6_lock : instruction_io_deq_ready_w_6_lock; // @[Decoder.scala 525:7 MultiEnqueue.scala 154:10]
  wire  _GEN_162 = _T_10 ? enqueuer4_io_in_ready : _GEN_124; // @[Decoder.scala 525:7 534:25]
  wire  _GEN_163 = _T_9 ? instruction_io_deq_valid : _GEN_125; // @[Decoder.scala 500:7 MultiEnqueue.scala 150:17]
  wire  _GEN_164 = _T_9 ? instruction_io_deq_ready_dataflow_io_enq_w_ready : _GEN_126; // @[Decoder.scala 500:7 ReadyValid.scala 19:11]
  wire  _GEN_165 = _T_9 ? instruction_io_deq_ready_dataflow_io_enq_w_2_valid : _GEN_127; // @[Decoder.scala 500:7 MultiEnqueue.scala 151:10]
  wire [3:0] _GEN_166 = _T_9 ? 4'h4 : _GEN_128; // @[Decoder.scala 500:7 MultiEnqueue.scala 151:10]
  wire [13:0] _GEN_167 = _T_9 ? instruction_io_deq_ready_w_size : _GEN_129; // @[Decoder.scala 500:7 MultiEnqueue.scala 151:10]
  wire  _GEN_168 = _T_9 ? instruction_io_deq_ready_lockPool_io_actor_0_in_w_ready : _GEN_130; // @[Decoder.scala 500:7 ReadyValid.scala 19:11]
  wire  _GEN_169 = _T_9 ? instruction_io_deq_ready_array_io_enq_w_3_valid : _GEN_131; // @[Decoder.scala 500:7 MultiEnqueue.scala 152:10]
  wire [13:0] _GEN_171 = _T_9 ? args_memAddress : _GEN_133; // @[Decoder.scala 500:7 MultiEnqueue.scala 152:10]
  wire [2:0] _GEN_173 = _T_9 ? args_memStride : _GEN_135; // @[Decoder.scala 500:7 MultiEnqueue.scala 152:10]
  wire  _GEN_175 = _T_9 ? instruction_io_deq_ready_acc_io_enq_w_ready : _GEN_137; // @[Decoder.scala 500:7 ReadyValid.scala 19:11]
  wire  _GEN_176 = _T_9 ? instruction_io_deq_ready_lockPool_io_actor_0_in_w_1_valid : _GEN_138; // @[Decoder.scala 500:7 MultiEnqueue.scala 153:10]
  wire [11:0] _GEN_181 = _T_9 ? instruction_io_deq_ready_w_2_address : _GEN_143; // @[Decoder.scala 500:7 MultiEnqueue.scala 153:10]
  wire  _GEN_184 = _T_9 ? 1'h0 : _GEN_146; // @[Decoder.scala 500:7 MultiEnqueue.scala 153:10]
  wire  _GEN_185 = _T_9 ? 1'h0 : _GEN_147; // @[Decoder.scala 500:7 MultiEnqueue.scala 153:10]
  wire [11:0] _GEN_186 = _T_9 ? instruction_io_deq_ready_w_2_size : _GEN_148; // @[Decoder.scala 500:7 MultiEnqueue.scala 153:10]
  wire [2:0] _GEN_187 = _T_9 ? args_accStride : _GEN_149; // @[Decoder.scala 500:7 MultiEnqueue.scala 153:10]
  wire  _GEN_189 = _T_9 ? instruction_io_deq_ready_lockPool_io_lock_w_ready : _GEN_151; // @[Decoder.scala 500:7 ReadyValid.scala 19:11]
  wire  _GEN_190 = _T_9 ? instruction_io_deq_ready_lockPool_io_lock_w_1_valid : _GEN_152; // @[Decoder.scala 500:7 MultiEnqueue.scala 154:10]
  wire [13:0] _GEN_193 = _T_9 ? instruction_io_deq_ready_w_size : _GEN_155; // @[Decoder.scala 500:7 MultiEnqueue.scala 154:10]
  wire  _GEN_196 = _T_9 ? instruction_io_deq_ready_w_6_lock : _GEN_158; // @[Decoder.scala 500:7 MultiEnqueue.scala 154:10]
  wire  _GEN_200 = _T_9 ? enqueuer4_io_in_ready : _GEN_162; // @[Decoder.scala 500:7 509:25]
  wire  _GEN_201 = _flags_WIRE_1 == 4'h3 ? instruction_io_deq_valid : _GEN_163; // @[Decoder.scala 470:59 MultiEnqueue.scala 150:17]
  wire  instruction_io_deq_ready_hostDataflow_io_enq_w_3_ready = hostDataflow_io_enq_ready; // @[MultiEnqueue.scala 151:10 ReadyValid.scala 16:17]
  wire  _GEN_202 = _flags_WIRE_1 == 4'h3 ? instruction_io_deq_ready_hostDataflow_io_enq_w_3_ready : _GEN_164; // @[Decoder.scala 470:59 ReadyValid.scala 19:11]
  wire  _GEN_203 = _flags_WIRE_1 == 4'h3 & instruction_io_deq_ready_dataflow_io_enq_w_2_valid; // @[Decoder.scala 470:59 MultiEnqueue.scala 151:10 Decoder.scala 670:16]
  wire [1:0] _GEN_204 = _flags_WIRE_1 == 4'h3 ? 2'h3 : 2'h0; // @[Decoder.scala 470:59 MultiEnqueue.scala 151:10 Decoder.scala 669:15]
  wire [13:0] _GEN_205 = _flags_WIRE_1 == 4'h3 ? instruction_io_deq_ready_w_size : 14'h0; // @[Decoder.scala 470:59 MultiEnqueue.scala 151:10 Decoder.scala 669:15]
  wire  instruction_io_deq_ready_lockPool_io_actor_1_in_w_3_ready = lockPool_io_actor_1_in_ready; // @[MultiEnqueue.scala 152:10 ReadyValid.scala 16:17]
  wire  _GEN_206 = _flags_WIRE_1 == 4'h3 ? instruction_io_deq_ready_lockPool_io_actor_1_in_w_3_ready : _GEN_168; // @[Decoder.scala 470:59 ReadyValid.scala 19:11]
  wire  _GEN_207 = _flags_WIRE_1 == 4'h3 & instruction_io_deq_ready_array_io_enq_w_3_valid; // @[Decoder.scala 470:59 MultiEnqueue.scala 152:10 Decoder.scala 670:16]
  wire [13:0] _GEN_209 = _flags_WIRE_1 == 4'h3 ? args_memAddress : 14'h0; // @[Decoder.scala 470:59 MultiEnqueue.scala 152:10 Decoder.scala 669:15]
  wire [2:0] _GEN_211 = _flags_WIRE_1 == 4'h3 ? args_memStride : 3'h0; // @[Decoder.scala 470:59 MultiEnqueue.scala 152:10 Decoder.scala 669:15]
  wire  instruction_io_deq_ready_dram1_io_enq_w_1_ready = dram1_io_enq_ready; // @[MultiEnqueue.scala 153:10 ReadyValid.scala 16:17]
  wire  _GEN_213 = _flags_WIRE_1 == 4'h3 ? instruction_io_deq_ready_dram1_io_enq_w_1_ready : _GEN_175; // @[Decoder.scala 470:59 ReadyValid.scala 19:11]
  wire  _GEN_214 = _flags_WIRE_1 == 4'h3 & instruction_io_deq_ready_lockPool_io_actor_0_in_w_1_valid; // @[Decoder.scala 470:59 MultiEnqueue.scala 153:10 Decoder.scala 670:16]
  wire [20:0] _GEN_216 = _flags_WIRE_1 == 4'h3 ? args_accAddress : 21'h0; // @[Decoder.scala 470:59 MultiEnqueue.scala 153:10 Decoder.scala 669:15]
  wire [20:0] instruction_io_deq_ready_w_21_size = {{5'd0}, args_size}; // @[MemControl.scala 44:19 46:14]
  wire [20:0] _GEN_217 = _flags_WIRE_1 == 4'h3 ? instruction_io_deq_ready_w_21_size : 21'h0; // @[Decoder.scala 470:59 MultiEnqueue.scala 153:10 Decoder.scala 669:15]
  wire [2:0] _GEN_218 = _flags_WIRE_1 == 4'h3 ? args_accStride : 3'h0; // @[Decoder.scala 470:59 MultiEnqueue.scala 153:10 Decoder.scala 669:15]
  wire  _GEN_220 = _flags_WIRE_1 == 4'h3 ? instruction_io_deq_ready_lockPool_io_lock_w_ready : _GEN_189; // @[Decoder.scala 470:59 ReadyValid.scala 19:11]
  wire  _GEN_221 = _flags_WIRE_1 == 4'h3 ? instruction_io_deq_ready_lockPool_io_lock_w_1_valid : _GEN_190; // @[Decoder.scala 470:59 MultiEnqueue.scala 154:10]
  wire  _GEN_222 = _flags_WIRE_1 == 4'h3 ? 1'h0 : _T_9; // @[Decoder.scala 470:59 MultiEnqueue.scala 154:10]
  wire [13:0] _GEN_224 = _flags_WIRE_1 == 4'h3 ? instruction_io_deq_ready_w_size : _GEN_193; // @[Decoder.scala 470:59 MultiEnqueue.scala 154:10]
  wire  _GEN_227 = _flags_WIRE_1 == 4'h3 ? instruction_io_deq_ready_w_6_lock : _GEN_196; // @[Decoder.scala 470:59 MultiEnqueue.scala 154:10]
  wire  _GEN_231 = _flags_WIRE_1 == 4'h3 ? enqueuer4_io_in_ready : _GEN_200; // @[Decoder.scala 470:59 478:25]
  wire  _GEN_232 = _flags_WIRE_1 == 4'h3 ? 1'h0 : _GEN_165; // @[Decoder.scala 470:59 670:16]
  wire [3:0] _GEN_233 = _flags_WIRE_1 == 4'h3 ? 4'h0 : _GEN_166; // @[Decoder.scala 470:59 669:15]
  wire [13:0] _GEN_234 = _flags_WIRE_1 == 4'h3 ? 14'h0 : _GEN_167; // @[Decoder.scala 470:59 669:15]
  wire  _GEN_235 = _flags_WIRE_1 == 4'h3 ? 1'h0 : _GEN_169; // @[Decoder.scala 470:59 670:16]
  wire [13:0] _GEN_237 = _flags_WIRE_1 == 4'h3 ? 14'h0 : _GEN_171; // @[Decoder.scala 470:59 669:15]
  wire [2:0] _GEN_239 = _flags_WIRE_1 == 4'h3 ? 3'h0 : _GEN_173; // @[Decoder.scala 470:59 669:15]
  wire  _GEN_241 = _flags_WIRE_1 == 4'h3 ? 1'h0 : _GEN_176; // @[Decoder.scala 470:59 670:16]
  wire [11:0] _GEN_246 = _flags_WIRE_1 == 4'h3 ? 12'h0 : _GEN_181; // @[Decoder.scala 470:59 669:15]
  wire  _GEN_249 = _flags_WIRE_1 == 4'h3 ? 1'h0 : _GEN_184; // @[Decoder.scala 470:59 669:15]
  wire  _GEN_250 = _flags_WIRE_1 == 4'h3 ? 1'h0 : _GEN_185; // @[Decoder.scala 470:59 669:15]
  wire [11:0] _GEN_251 = _flags_WIRE_1 == 4'h3 ? 12'h0 : _GEN_186; // @[Decoder.scala 470:59 669:15]
  wire [2:0] _GEN_252 = _flags_WIRE_1 == 4'h3 ? 3'h0 : _GEN_187; // @[Decoder.scala 470:59 669:15]
  wire  _GEN_254 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_valid : _GEN_201; // @[Decoder.scala 441:59 MultiEnqueue.scala 150:17]
  wire  _GEN_255 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_hostDataflow_io_enq_w_3_ready : _GEN_202; // @[Decoder.scala 441:59 ReadyValid.scala 19:11]
  wire  _GEN_256 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_dataflow_io_enq_w_2_valid : _GEN_203; // @[Decoder.scala 441:59 MultiEnqueue.scala 151:10]
  wire [1:0] _GEN_257 = _flags_WIRE_1 == 4'h2 ? 2'h2 : _GEN_204; // @[Decoder.scala 441:59 MultiEnqueue.scala 151:10]
  wire [13:0] _GEN_258 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_w_size : _GEN_205; // @[Decoder.scala 441:59 MultiEnqueue.scala 151:10]
  wire  _GEN_259 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_lockPool_io_actor_1_in_w_3_ready : _GEN_206; // @[Decoder.scala 441:59 ReadyValid.scala 19:11]
  wire  _GEN_260 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_array_io_enq_w_3_valid : _GEN_207; // @[Decoder.scala 441:59 MultiEnqueue.scala 152:10]
  wire [13:0] _GEN_262 = _flags_WIRE_1 == 4'h2 ? args_memAddress : _GEN_209; // @[Decoder.scala 441:59 MultiEnqueue.scala 152:10]
  wire [2:0] _GEN_264 = _flags_WIRE_1 == 4'h2 ? args_memStride : _GEN_211; // @[Decoder.scala 441:59 MultiEnqueue.scala 152:10]
  wire  _GEN_266 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_dram1_io_enq_w_1_ready : _GEN_213; // @[Decoder.scala 441:59 ReadyValid.scala 19:11]
  wire  _GEN_267 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_lockPool_io_actor_0_in_w_1_valid : _GEN_214; // @[Decoder.scala 441:59 MultiEnqueue.scala 153:10]
  wire  _GEN_268 = _flags_WIRE_1 == 4'h2 ? 1'h0 : _T_8; // @[Decoder.scala 441:59 MultiEnqueue.scala 153:10]
  wire [20:0] _GEN_269 = _flags_WIRE_1 == 4'h2 ? args_accAddress : _GEN_216; // @[Decoder.scala 441:59 MultiEnqueue.scala 153:10]
  wire [20:0] _GEN_270 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_w_21_size : _GEN_217; // @[Decoder.scala 441:59 MultiEnqueue.scala 153:10]
  wire [2:0] _GEN_271 = _flags_WIRE_1 == 4'h2 ? args_accStride : _GEN_218; // @[Decoder.scala 441:59 MultiEnqueue.scala 153:10]
  wire  _GEN_273 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_lockPool_io_lock_w_ready : _GEN_220; // @[Decoder.scala 441:59 ReadyValid.scala 19:11]
  wire  _GEN_274 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_lockPool_io_lock_w_1_valid : _GEN_221; // @[Decoder.scala 441:59 MultiEnqueue.scala 154:10]
  wire  _GEN_275 = _flags_WIRE_1 == 4'h2 | _GEN_222; // @[Decoder.scala 441:59 MultiEnqueue.scala 154:10]
  wire [13:0] _GEN_277 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_w_size : _GEN_224; // @[Decoder.scala 441:59 MultiEnqueue.scala 154:10]
  wire  _GEN_280 = _flags_WIRE_1 == 4'h2 ? instruction_io_deq_ready_w_6_lock : _GEN_227; // @[Decoder.scala 441:59 MultiEnqueue.scala 154:10]
  wire  _GEN_282 = _flags_WIRE_1 == 4'h2 | _T_8; // @[Decoder.scala 441:59 MultiEnqueue.scala 154:10]
  wire  _GEN_284 = _flags_WIRE_1 == 4'h2 ? enqueuer4_io_in_ready : _GEN_231; // @[Decoder.scala 441:59 450:25]
  wire  _GEN_285 = _flags_WIRE_1 == 4'h2 ? 1'h0 : _GEN_232; // @[Decoder.scala 441:59 670:16]
  wire [3:0] _GEN_286 = _flags_WIRE_1 == 4'h2 ? 4'h0 : _GEN_233; // @[Decoder.scala 441:59 669:15]
  wire [13:0] _GEN_287 = _flags_WIRE_1 == 4'h2 ? 14'h0 : _GEN_234; // @[Decoder.scala 441:59 669:15]
  wire  _GEN_288 = _flags_WIRE_1 == 4'h2 ? 1'h0 : _GEN_235; // @[Decoder.scala 441:59 670:16]
  wire  _GEN_289 = _flags_WIRE_1 == 4'h2 ? 1'h0 : _GEN_222; // @[Decoder.scala 441:59 669:15]
  wire [13:0] _GEN_290 = _flags_WIRE_1 == 4'h2 ? 14'h0 : _GEN_237; // @[Decoder.scala 441:59 669:15]
  wire [2:0] _GEN_292 = _flags_WIRE_1 == 4'h2 ? 3'h0 : _GEN_239; // @[Decoder.scala 441:59 669:15]
  wire  _GEN_294 = _flags_WIRE_1 == 4'h2 ? 1'h0 : _GEN_241; // @[Decoder.scala 441:59 670:16]
  wire [11:0] _GEN_299 = _flags_WIRE_1 == 4'h2 ? 12'h0 : _GEN_246; // @[Decoder.scala 441:59 669:15]
  wire  _GEN_302 = _flags_WIRE_1 == 4'h2 ? 1'h0 : _GEN_249; // @[Decoder.scala 441:59 669:15]
  wire  _GEN_303 = _flags_WIRE_1 == 4'h2 ? 1'h0 : _GEN_250; // @[Decoder.scala 441:59 669:15]
  wire [11:0] _GEN_304 = _flags_WIRE_1 == 4'h2 ? 12'h0 : _GEN_251; // @[Decoder.scala 441:59 669:15]
  wire [2:0] _GEN_305 = _flags_WIRE_1 == 4'h2 ? 3'h0 : _GEN_252; // @[Decoder.scala 441:59 669:15]
  wire  _GEN_307 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_valid : _GEN_254; // @[Decoder.scala 412:59 MultiEnqueue.scala 150:17]
  wire  _GEN_308 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_hostDataflow_io_enq_w_3_ready : _GEN_255; // @[Decoder.scala 412:59 ReadyValid.scala 19:11]
  wire  _GEN_309 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_dataflow_io_enq_w_2_valid : _GEN_256; // @[Decoder.scala 412:59 MultiEnqueue.scala 151:10]
  wire [1:0] _GEN_310 = _flags_WIRE_1 == 4'h1 ? 2'h1 : _GEN_257; // @[Decoder.scala 412:59 MultiEnqueue.scala 151:10]
  wire [13:0] _GEN_311 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_w_size : _GEN_258; // @[Decoder.scala 412:59 MultiEnqueue.scala 151:10]
  wire  _GEN_312 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_lockPool_io_actor_1_in_w_3_ready : _GEN_259; // @[Decoder.scala 412:59 ReadyValid.scala 19:11]
  wire  _GEN_313 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_array_io_enq_w_3_valid : _GEN_260; // @[Decoder.scala 412:59 MultiEnqueue.scala 152:10]
  wire  _GEN_314 = _flags_WIRE_1 == 4'h1 ? 1'h0 : _T_7; // @[Decoder.scala 412:59 MultiEnqueue.scala 152:10]
  wire [13:0] _GEN_315 = _flags_WIRE_1 == 4'h1 ? args_memAddress : _GEN_262; // @[Decoder.scala 412:59 MultiEnqueue.scala 152:10]
  wire [2:0] _GEN_317 = _flags_WIRE_1 == 4'h1 ? args_memStride : _GEN_264; // @[Decoder.scala 412:59 MultiEnqueue.scala 152:10]
  wire  instruction_io_deq_ready_dram0_io_enq_w_1_ready = dram0_io_enq_ready; // @[MultiEnqueue.scala 153:10 ReadyValid.scala 16:17]
  wire  _GEN_319 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_dram0_io_enq_w_1_ready : _GEN_266; // @[Decoder.scala 412:59 ReadyValid.scala 19:11]
  wire  _GEN_320 = _flags_WIRE_1 == 4'h1 & instruction_io_deq_ready_lockPool_io_actor_0_in_w_1_valid; // @[Decoder.scala 412:59 MultiEnqueue.scala 153:10 Decoder.scala 670:16]
  wire [20:0] _GEN_322 = _flags_WIRE_1 == 4'h1 ? args_accAddress : 21'h0; // @[Decoder.scala 412:59 MultiEnqueue.scala 153:10 Decoder.scala 669:15]
  wire [20:0] _GEN_323 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_w_21_size : 21'h0; // @[Decoder.scala 412:59 MultiEnqueue.scala 153:10 Decoder.scala 669:15]
  wire [2:0] _GEN_324 = _flags_WIRE_1 == 4'h1 ? args_accStride : 3'h0; // @[Decoder.scala 412:59 MultiEnqueue.scala 153:10 Decoder.scala 669:15]
  wire  _GEN_326 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_lockPool_io_lock_w_ready : _GEN_273; // @[Decoder.scala 412:59 ReadyValid.scala 19:11]
  wire  _GEN_327 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_lockPool_io_lock_w_1_valid : _GEN_274; // @[Decoder.scala 412:59 MultiEnqueue.scala 154:10]
  wire  _GEN_328 = _flags_WIRE_1 == 4'h1 ? 1'h0 : _GEN_275; // @[Decoder.scala 412:59 MultiEnqueue.scala 154:10]
  wire [13:0] _GEN_330 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_w_size : _GEN_277; // @[Decoder.scala 412:59 MultiEnqueue.scala 154:10]
  wire  _GEN_333 = _flags_WIRE_1 == 4'h1 ? instruction_io_deq_ready_w_6_lock : _GEN_280; // @[Decoder.scala 412:59 MultiEnqueue.scala 154:10]
  wire  _GEN_335 = _flags_WIRE_1 == 4'h1 | _GEN_282; // @[Decoder.scala 412:59 MultiEnqueue.scala 154:10]
  wire  _GEN_337 = _flags_WIRE_1 == 4'h1 ? enqueuer4_io_in_ready : _GEN_284; // @[Decoder.scala 412:59 421:25]
  wire  _GEN_338 = _flags_WIRE_1 == 4'h1 ? 1'h0 : _GEN_267; // @[Decoder.scala 412:59 670:16]
  wire  _GEN_339 = _flags_WIRE_1 == 4'h1 ? 1'h0 : _GEN_268; // @[Decoder.scala 412:59 669:15]
  wire [20:0] _GEN_340 = _flags_WIRE_1 == 4'h1 ? 21'h0 : _GEN_269; // @[Decoder.scala 412:59 669:15]
  wire [20:0] _GEN_341 = _flags_WIRE_1 == 4'h1 ? 21'h0 : _GEN_270; // @[Decoder.scala 412:59 669:15]
  wire [2:0] _GEN_342 = _flags_WIRE_1 == 4'h1 ? 3'h0 : _GEN_271; // @[Decoder.scala 412:59 669:15]
  wire  _GEN_344 = _flags_WIRE_1 == 4'h1 ? 1'h0 : _GEN_285; // @[Decoder.scala 412:59 670:16]
  wire [3:0] _GEN_345 = _flags_WIRE_1 == 4'h1 ? 4'h0 : _GEN_286; // @[Decoder.scala 412:59 669:15]
  wire [13:0] _GEN_346 = _flags_WIRE_1 == 4'h1 ? 14'h0 : _GEN_287; // @[Decoder.scala 412:59 669:15]
  wire  _GEN_347 = _flags_WIRE_1 == 4'h1 ? 1'h0 : _GEN_288; // @[Decoder.scala 412:59 670:16]
  wire  _GEN_348 = _flags_WIRE_1 == 4'h1 ? 1'h0 : _GEN_289; // @[Decoder.scala 412:59 669:15]
  wire [13:0] _GEN_349 = _flags_WIRE_1 == 4'h1 ? 14'h0 : _GEN_290; // @[Decoder.scala 412:59 669:15]
  wire [2:0] _GEN_351 = _flags_WIRE_1 == 4'h1 ? 3'h0 : _GEN_292; // @[Decoder.scala 412:59 669:15]
  wire  _GEN_353 = _flags_WIRE_1 == 4'h1 ? 1'h0 : _GEN_294; // @[Decoder.scala 412:59 670:16]
  wire [11:0] _GEN_358 = _flags_WIRE_1 == 4'h1 ? 12'h0 : _GEN_299; // @[Decoder.scala 412:59 669:15]
  wire  _GEN_361 = _flags_WIRE_1 == 4'h1 ? 1'h0 : _GEN_302; // @[Decoder.scala 412:59 669:15]
  wire  _GEN_362 = _flags_WIRE_1 == 4'h1 ? 1'h0 : _GEN_303; // @[Decoder.scala 412:59 669:15]
  wire [11:0] _GEN_363 = _flags_WIRE_1 == 4'h1 ? 12'h0 : _GEN_304; // @[Decoder.scala 412:59 669:15]
  wire [2:0] _GEN_364 = _flags_WIRE_1 == 4'h1 ? 3'h0 : _GEN_305; // @[Decoder.scala 412:59 669:15]
  wire  _GEN_366 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_valid : _GEN_307; // @[Decoder.scala 383:53 MultiEnqueue.scala 150:17]
  wire  _GEN_367 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_hostDataflow_io_enq_w_3_ready : _GEN_308; // @[Decoder.scala 383:53 ReadyValid.scala 19:11]
  wire  _GEN_368 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_dataflow_io_enq_w_2_valid : _GEN_309; // @[Decoder.scala 383:53 MultiEnqueue.scala 151:10]
  wire [1:0] _GEN_369 = _flags_WIRE_1 == 4'h0 ? 2'h0 : _GEN_310; // @[Decoder.scala 383:53 MultiEnqueue.scala 151:10]
  wire [13:0] _GEN_370 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_w_size : _GEN_311; // @[Decoder.scala 383:53 MultiEnqueue.scala 151:10]
  wire  _GEN_371 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_lockPool_io_actor_1_in_w_3_ready : _GEN_312; // @[Decoder.scala 383:53 ReadyValid.scala 19:11]
  wire  _GEN_372 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_array_io_enq_w_3_valid : _GEN_313; // @[Decoder.scala 383:53 MultiEnqueue.scala 152:10]
  wire  _GEN_373 = _flags_WIRE_1 == 4'h0 | _GEN_314; // @[Decoder.scala 383:53 MultiEnqueue.scala 152:10]
  wire [13:0] _GEN_374 = _flags_WIRE_1 == 4'h0 ? args_memAddress : _GEN_315; // @[Decoder.scala 383:53 MultiEnqueue.scala 152:10]
  wire [2:0] _GEN_376 = _flags_WIRE_1 == 4'h0 ? args_memStride : _GEN_317; // @[Decoder.scala 383:53 MultiEnqueue.scala 152:10]
  wire  _GEN_378 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_dram0_io_enq_w_1_ready : _GEN_319; // @[Decoder.scala 383:53 ReadyValid.scala 19:11]
  wire  _GEN_379 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_lockPool_io_actor_0_in_w_1_valid : _GEN_320; // @[Decoder.scala 383:53 MultiEnqueue.scala 153:10]
  wire  _GEN_380 = _flags_WIRE_1 == 4'h0 ? 1'h0 : _T_6; // @[Decoder.scala 383:53 MultiEnqueue.scala 153:10]
  wire [20:0] _GEN_381 = _flags_WIRE_1 == 4'h0 ? args_accAddress : _GEN_322; // @[Decoder.scala 383:53 MultiEnqueue.scala 153:10]
  wire [20:0] _GEN_382 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_w_21_size : _GEN_323; // @[Decoder.scala 383:53 MultiEnqueue.scala 153:10]
  wire [2:0] _GEN_383 = _flags_WIRE_1 == 4'h0 ? args_accStride : _GEN_324; // @[Decoder.scala 383:53 MultiEnqueue.scala 153:10]
  wire  _GEN_385 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_lockPool_io_lock_w_ready : _GEN_326; // @[Decoder.scala 383:53 ReadyValid.scala 19:11]
  wire  _GEN_386 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_lockPool_io_lock_w_1_valid : _GEN_327; // @[Decoder.scala 383:53 MultiEnqueue.scala 154:10]
  wire  _GEN_387 = _flags_WIRE_1 == 4'h0 | _GEN_328; // @[Decoder.scala 383:53 MultiEnqueue.scala 154:10]
  wire [13:0] _GEN_389 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_w_size : _GEN_330; // @[Decoder.scala 383:53 MultiEnqueue.scala 154:10]
  wire  _GEN_392 = _flags_WIRE_1 == 4'h0 ? instruction_io_deq_ready_w_6_lock : _GEN_333; // @[Decoder.scala 383:53 MultiEnqueue.scala 154:10]
  wire  _GEN_394 = _flags_WIRE_1 == 4'h0 | _GEN_335; // @[Decoder.scala 383:53 MultiEnqueue.scala 154:10]
  wire  _GEN_396 = _flags_WIRE_1 == 4'h0 ? enqueuer4_io_in_ready : _GEN_337; // @[Decoder.scala 383:53 392:25]
  wire  _GEN_397 = _flags_WIRE_1 == 4'h0 ? 1'h0 : _GEN_338; // @[Decoder.scala 383:53 670:16]
  wire  _GEN_398 = _flags_WIRE_1 == 4'h0 ? 1'h0 : _GEN_339; // @[Decoder.scala 383:53 669:15]
  wire [20:0] _GEN_399 = _flags_WIRE_1 == 4'h0 ? 21'h0 : _GEN_340; // @[Decoder.scala 383:53 669:15]
  wire [20:0] _GEN_400 = _flags_WIRE_1 == 4'h0 ? 21'h0 : _GEN_341; // @[Decoder.scala 383:53 669:15]
  wire [2:0] _GEN_401 = _flags_WIRE_1 == 4'h0 ? 3'h0 : _GEN_342; // @[Decoder.scala 383:53 669:15]
  wire  _GEN_403 = _flags_WIRE_1 == 4'h0 ? 1'h0 : _GEN_344; // @[Decoder.scala 383:53 670:16]
  wire [3:0] _GEN_404 = _flags_WIRE_1 == 4'h0 ? 4'h0 : _GEN_345; // @[Decoder.scala 383:53 669:15]
  wire [13:0] _GEN_405 = _flags_WIRE_1 == 4'h0 ? 14'h0 : _GEN_346; // @[Decoder.scala 383:53 669:15]
  wire  _GEN_406 = _flags_WIRE_1 == 4'h0 ? 1'h0 : _GEN_347; // @[Decoder.scala 383:53 670:16]
  wire  _GEN_407 = _flags_WIRE_1 == 4'h0 ? 1'h0 : _GEN_348; // @[Decoder.scala 383:53 669:15]
  wire [13:0] _GEN_408 = _flags_WIRE_1 == 4'h0 ? 14'h0 : _GEN_349; // @[Decoder.scala 383:53 669:15]
  wire [2:0] _GEN_410 = _flags_WIRE_1 == 4'h0 ? 3'h0 : _GEN_351; // @[Decoder.scala 383:53 669:15]
  wire  _GEN_412 = _flags_WIRE_1 == 4'h0 ? 1'h0 : _GEN_353; // @[Decoder.scala 383:53 670:16]
  wire [11:0] _GEN_417 = _flags_WIRE_1 == 4'h0 ? 12'h0 : _GEN_358; // @[Decoder.scala 383:53 669:15]
  wire  _GEN_420 = _flags_WIRE_1 == 4'h0 ? 1'h0 : _GEN_361; // @[Decoder.scala 383:53 669:15]
  wire  _GEN_421 = _flags_WIRE_1 == 4'h0 ? 1'h0 : _GEN_362; // @[Decoder.scala 383:53 669:15]
  wire [11:0] _GEN_422 = _flags_WIRE_1 == 4'h0 ? 12'h0 : _GEN_363; // @[Decoder.scala 383:53 669:15]
  wire [2:0] _GEN_423 = _flags_WIRE_1 == 4'h0 ? 3'h0 : _GEN_364; // @[Decoder.scala 383:53 669:15]
  wire  flags_3_accumulate = _flags_WIRE_1[2]; // @[Decoder.scala 583:45]
  wire [23:0] args_3_accWriteAddress = _args_WIRE_1[23:0]; // @[Decoder.scala 584:48]
  wire [23:0] args_3_accReadAddress = _args_WIRE_1[47:24]; // @[Decoder.scala 584:48]
  wire  args_3_instruction_dest = _args_WIRE_1[48]; // @[Decoder.scala 584:48]
  wire  args_3_instruction_sourceRight = _args_WIRE_1[49]; // @[Decoder.scala 584:48]
  wire  args_3_instruction_sourceLeft = _args_WIRE_1[50]; // @[Decoder.scala 584:48]
  wire [3:0] args_3_instruction_op = _args_WIRE_1[54:51]; // @[Decoder.scala 584:48]
  wire [3:0] args_4_register = instruction_io_deq_bits_arguments[3:0]; // @[Decoder.scala 610:50]
  wire [27:0] args_4_value = instruction_io_deq_bits_arguments[31:4]; // @[Decoder.scala 610:50]
  wire [43:0] _dram0AddressOffset_T = {args_4_value, 16'h0}; // @[Decoder.scala 613:43]
  wire [31:0] _GEN_426 = args_4_register == 4'ha ? {{4'd0}, args_4_value} : _GEN_2; // @[Decoder.scala 624:62 625:24]
  wire [31:0] _GEN_428 = args_4_register == 4'h9 ? {{4'd0}, args_4_value} : tracepoint; // @[Decoder.scala 622:58 623:20 108:31]
  wire [31:0] _GEN_429 = args_4_register == 4'h9 ? _GEN_2 : _GEN_426; // @[Decoder.scala 622:58]
  wire [27:0] _GEN_431 = args_4_register == 4'h8 ? args_4_value : {{12'd0}, timeout}; // @[Decoder.scala 620:55 621:17 96:24]
  wire [31:0] _GEN_432 = args_4_register == 4'h8 ? tracepoint : _GEN_428; // @[Decoder.scala 108:31 620:55]
  wire [31:0] _GEN_433 = args_4_register == 4'h8 ? _GEN_2 : _GEN_429; // @[Decoder.scala 620:55]
  wire [27:0] _GEN_435 = args_4_register == 4'h5 ? args_4_value : {{24'd0}, dram1CacheBehaviour}; // @[Decoder.scala 618:67 619:29 133:36]
  wire [27:0] _GEN_436 = args_4_register == 4'h5 ? {{12'd0}, timeout} : _GEN_431; // @[Decoder.scala 618:67 96:24]
  wire [31:0] _GEN_437 = args_4_register == 4'h5 ? tracepoint : _GEN_432; // @[Decoder.scala 108:31 618:67]
  wire [31:0] _GEN_438 = args_4_register == 4'h5 ? _GEN_2 : _GEN_433; // @[Decoder.scala 618:67]
  wire [43:0] _GEN_440 = args_4_register == 4'h4 ? _dram0AddressOffset_T : {{12'd0}, dram1AddressOffset}; // @[Decoder.scala 616:66 617:28 130:35]
  wire [27:0] _GEN_441 = args_4_register == 4'h4 ? {{24'd0}, dram1CacheBehaviour} : _GEN_435; // @[Decoder.scala 133:36 616:66]
  wire [27:0] _GEN_442 = args_4_register == 4'h4 ? {{12'd0}, timeout} : _GEN_436; // @[Decoder.scala 616:66 96:24]
  wire [31:0] _GEN_443 = args_4_register == 4'h4 ? tracepoint : _GEN_437; // @[Decoder.scala 108:31 616:66]
  wire [31:0] _GEN_444 = args_4_register == 4'h4 ? _GEN_2 : _GEN_438; // @[Decoder.scala 616:66]
  wire [27:0] _GEN_446 = args_4_register == 4'h1 ? args_4_value : {{24'd0}, dram0CacheBehaviour}; // @[Decoder.scala 614:67 615:29 129:36]
  wire [43:0] _GEN_447 = args_4_register == 4'h1 ? {{12'd0}, dram1AddressOffset} : _GEN_440; // @[Decoder.scala 130:35 614:67]
  wire [27:0] _GEN_448 = args_4_register == 4'h1 ? {{24'd0}, dram1CacheBehaviour} : _GEN_441; // @[Decoder.scala 133:36 614:67]
  wire [27:0] _GEN_449 = args_4_register == 4'h1 ? {{12'd0}, timeout} : _GEN_442; // @[Decoder.scala 614:67 96:24]
  wire [31:0] _GEN_450 = args_4_register == 4'h1 ? tracepoint : _GEN_443; // @[Decoder.scala 108:31 614:67]
  wire [31:0] _GEN_451 = args_4_register == 4'h1 ? _GEN_2 : _GEN_444; // @[Decoder.scala 614:67]
  wire [43:0] _GEN_453 = args_4_register == 4'h0 ? _dram0AddressOffset_T : {{12'd0}, dram0AddressOffset}; // @[Decoder.scala 612:60 613:28 126:35]
  wire [27:0] _GEN_454 = args_4_register == 4'h0 ? {{24'd0}, dram0CacheBehaviour} : _GEN_446; // @[Decoder.scala 129:36 612:60]
  wire [43:0] _GEN_455 = args_4_register == 4'h0 ? {{12'd0}, dram1AddressOffset} : _GEN_447; // @[Decoder.scala 130:35 612:60]
  wire [27:0] _GEN_456 = args_4_register == 4'h0 ? {{24'd0}, dram1CacheBehaviour} : _GEN_448; // @[Decoder.scala 133:36 612:60]
  wire [27:0] _GEN_457 = args_4_register == 4'h0 ? {{12'd0}, timeout} : _GEN_449; // @[Decoder.scala 612:60 96:24]
  wire [31:0] _GEN_458 = args_4_register == 4'h0 ? tracepoint : _GEN_450; // @[Decoder.scala 108:31 612:60]
  wire [31:0] _GEN_459 = args_4_register == 4'h0 ? _GEN_2 : _GEN_451; // @[Decoder.scala 612:60]
  wire [43:0] _GEN_461 = instruction_io_deq_valid ? _GEN_453 : {{12'd0}, dram0AddressOffset}; // @[Decoder.scala 601:29 126:35]
  wire [27:0] _GEN_462 = instruction_io_deq_valid ? _GEN_454 : {{24'd0}, dram0CacheBehaviour}; // @[Decoder.scala 601:29 129:36]
  wire [43:0] _GEN_463 = instruction_io_deq_valid ? _GEN_455 : {{12'd0}, dram1AddressOffset}; // @[Decoder.scala 601:29 130:35]
  wire [27:0] _GEN_464 = instruction_io_deq_valid ? _GEN_456 : {{24'd0}, dram1CacheBehaviour}; // @[Decoder.scala 601:29 133:36]
  wire [27:0] _GEN_465 = instruction_io_deq_valid ? _GEN_457 : {{12'd0}, timeout}; // @[Decoder.scala 601:29 96:24]
  wire [31:0] _GEN_466 = instruction_io_deq_valid ? _GEN_458 : tracepoint; // @[Decoder.scala 601:29 108:31]
  wire [31:0] _GEN_467 = instruction_io_deq_valid ? _GEN_459 : _GEN_2; // @[Decoder.scala 601:29]
  wire [43:0] _GEN_472 = instruction_io_deq_bits_opcode == 4'hf ? _GEN_461 : {{12'd0}, dram0AddressOffset}; // @[Decoder.scala 126:35 600:60]
  wire [27:0] _GEN_473 = instruction_io_deq_bits_opcode == 4'hf ? _GEN_462 : {{24'd0}, dram0CacheBehaviour}; // @[Decoder.scala 129:36 600:60]
  wire [43:0] _GEN_474 = instruction_io_deq_bits_opcode == 4'hf ? _GEN_463 : {{12'd0}, dram1AddressOffset}; // @[Decoder.scala 130:35 600:60]
  wire [27:0] _GEN_475 = instruction_io_deq_bits_opcode == 4'hf ? _GEN_464 : {{24'd0}, dram1CacheBehaviour}; // @[Decoder.scala 133:36 600:60]
  wire [27:0] _GEN_476 = instruction_io_deq_bits_opcode == 4'hf ? _GEN_465 : {{12'd0}, timeout}; // @[Decoder.scala 600:60 96:24]
  wire [31:0] _GEN_477 = instruction_io_deq_bits_opcode == 4'hf ? _GEN_466 : tracepoint; // @[Decoder.scala 108:31 600:60]
  wire [31:0] _GEN_478 = instruction_io_deq_bits_opcode == 4'hf ? _GEN_467 : _GEN_2; // @[Decoder.scala 600:60]
  wire  _GEN_483 = instruction_io_deq_bits_opcode == 4'h4 & instruction_io_deq_valid; // @[Decoder.scala 577:55 MultiEnqueue.scala 40:17 60:17]
  wire  _GEN_484 = instruction_io_deq_bits_opcode == 4'h4 & instruction_io_deq_ready_acc_io_enq_w_ready; // @[Decoder.scala 577:55 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  _GEN_485 = instruction_io_deq_bits_opcode == 4'h4 & instruction_io_deq_ready_array_io_enq_w_2_valid; // @[Decoder.scala 577:55 MultiEnqueue.scala 61:10 Decoder.scala 670:16]
  wire [3:0] _GEN_486 = instruction_io_deq_bits_opcode == 4'h4 ? args_3_instruction_op : 4'h0; // @[Decoder.scala 577:55 MultiEnqueue.scala 61:10 Decoder.scala 669:15]
  wire  _GEN_487 = instruction_io_deq_bits_opcode == 4'h4 & args_3_instruction_sourceLeft; // @[Decoder.scala 577:55 MultiEnqueue.scala 61:10 Decoder.scala 669:15]
  wire  _GEN_488 = instruction_io_deq_bits_opcode == 4'h4 & args_3_instruction_sourceRight; // @[Decoder.scala 577:55 MultiEnqueue.scala 61:10 Decoder.scala 669:15]
  wire  _GEN_489 = instruction_io_deq_bits_opcode == 4'h4 & args_3_instruction_dest; // @[Decoder.scala 577:55 MultiEnqueue.scala 61:10 Decoder.scala 669:15]
  wire [11:0] instruction_io_deq_ready_w_32_address = args_3_accReadAddress[11:0]; // @[Decoder.scala 716:17 718:15]
  wire [11:0] _GEN_490 = instruction_io_deq_bits_opcode == 4'h4 ? instruction_io_deq_ready_w_32_address : 12'h0; // @[Decoder.scala 577:55 MultiEnqueue.scala 61:10 Decoder.scala 669:15]
  wire [11:0] instruction_io_deq_ready_w_32_altAddress = args_3_accWriteAddress[11:0]; // @[Decoder.scala 716:17 719:18]
  wire [11:0] _GEN_491 = instruction_io_deq_bits_opcode == 4'h4 ? instruction_io_deq_ready_w_32_altAddress : 12'h0; // @[Decoder.scala 577:55 MultiEnqueue.scala 61:10 Decoder.scala 669:15]
  wire  _GEN_492 = instruction_io_deq_bits_opcode == 4'h4 & flags_accumulate; // @[Decoder.scala 577:55 MultiEnqueue.scala 61:10 Decoder.scala 669:15]
  wire  _GEN_493 = instruction_io_deq_bits_opcode == 4'h4 & flags_zeroes; // @[Decoder.scala 577:55 MultiEnqueue.scala 61:10 Decoder.scala 669:15]
  wire  _GEN_494 = instruction_io_deq_bits_opcode == 4'h4 & flags_3_accumulate; // @[Decoder.scala 577:55 MultiEnqueue.scala 61:10 Decoder.scala 669:15]
  wire  _GEN_498 = instruction_io_deq_bits_opcode == 4'h4 ? enqueuer1_io_in_ready : 1'h1; // @[Decoder.scala 577:55 586:23]
  wire [43:0] _GEN_499 = instruction_io_deq_bits_opcode == 4'h4 ? {{12'd0}, dram0AddressOffset} : _GEN_472; // @[Decoder.scala 126:35 577:55]
  wire [27:0] _GEN_500 = instruction_io_deq_bits_opcode == 4'h4 ? {{24'd0}, dram0CacheBehaviour} : _GEN_473; // @[Decoder.scala 129:36 577:55]
  wire [43:0] _GEN_501 = instruction_io_deq_bits_opcode == 4'h4 ? {{12'd0}, dram1AddressOffset} : _GEN_474; // @[Decoder.scala 130:35 577:55]
  wire [27:0] _GEN_502 = instruction_io_deq_bits_opcode == 4'h4 ? {{24'd0}, dram1CacheBehaviour} : _GEN_475; // @[Decoder.scala 133:36 577:55]
  wire [27:0] _GEN_503 = instruction_io_deq_bits_opcode == 4'h4 ? {{12'd0}, timeout} : _GEN_476; // @[Decoder.scala 577:55 96:24]
  wire [31:0] _GEN_504 = instruction_io_deq_bits_opcode == 4'h4 ? tracepoint : _GEN_477; // @[Decoder.scala 108:31 577:55]
  wire [31:0] _GEN_505 = instruction_io_deq_bits_opcode == 4'h4 ? _GEN_2 : _GEN_478; // @[Decoder.scala 577:55]
  wire  _GEN_509 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_366; // @[Decoder.scala 373:59 MultiEnqueue.scala 40:17]
  wire  _GEN_510 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_367; // @[Decoder.scala 373:59 MultiEnqueue.scala 42:18]
  wire  _GEN_511 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_368; // @[Decoder.scala 373:59 670:16]
  wire [1:0] _GEN_512 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_369 : 2'h0; // @[Decoder.scala 373:59 669:15]
  wire [13:0] _GEN_513 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_370 : 14'h0; // @[Decoder.scala 373:59 669:15]
  wire  _GEN_514 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_371; // @[Decoder.scala 373:59 MultiEnqueue.scala 42:18]
  wire  _GEN_515 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_372; // @[Decoder.scala 373:59 670:16]
  wire  _GEN_516 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_373; // @[Decoder.scala 373:59 669:15]
  wire [13:0] _GEN_517 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_374 : 14'h0; // @[Decoder.scala 373:59 669:15]
  wire [2:0] _GEN_519 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_376 : 3'h0; // @[Decoder.scala 373:59 669:15]
  wire  _GEN_521 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_378; // @[Decoder.scala 373:59 MultiEnqueue.scala 42:18]
  wire  _GEN_522 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_379; // @[Decoder.scala 373:59 670:16]
  wire  _GEN_523 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_380; // @[Decoder.scala 373:59 669:15]
  wire [20:0] _GEN_524 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_381 : 21'h0; // @[Decoder.scala 373:59 669:15]
  wire [20:0] _GEN_525 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_382 : 21'h0; // @[Decoder.scala 373:59 669:15]
  wire [2:0] _GEN_526 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_383 : 3'h0; // @[Decoder.scala 373:59 669:15]
  wire  _GEN_528 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_385; // @[Decoder.scala 373:59 MultiEnqueue.scala 42:18]
  wire  _GEN_529 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_386; // @[Decoder.scala 373:59 Decoupled.scala 72:20]
  wire  _GEN_539 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_396 : _GEN_498; // @[Decoder.scala 373:59]
  wire  _GEN_540 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_397; // @[Decoder.scala 373:59 670:16]
  wire  _GEN_541 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_398; // @[Decoder.scala 373:59 669:15]
  wire [20:0] _GEN_542 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_399 : 21'h0; // @[Decoder.scala 373:59 669:15]
  wire [20:0] _GEN_543 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_400 : 21'h0; // @[Decoder.scala 373:59 669:15]
  wire [2:0] _GEN_544 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_401 : 3'h0; // @[Decoder.scala 373:59 669:15]
  wire  _GEN_546 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_403; // @[Decoder.scala 373:59 670:16]
  wire [3:0] _GEN_547 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_404 : 4'h0; // @[Decoder.scala 373:59 669:15]
  wire [13:0] _GEN_548 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_405 : 14'h0; // @[Decoder.scala 373:59 669:15]
  wire  _GEN_549 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_406; // @[Decoder.scala 373:59 670:16]
  wire  _GEN_550 = instruction_io_deq_bits_opcode == 4'h2 & _GEN_407; // @[Decoder.scala 373:59 669:15]
  wire [13:0] _GEN_551 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_408 : 14'h0; // @[Decoder.scala 373:59 669:15]
  wire [2:0] _GEN_553 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_410 : 3'h0; // @[Decoder.scala 373:59 669:15]
  wire  _GEN_555 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_412 : _GEN_485; // @[Decoder.scala 373:59]
  wire [3:0] _GEN_556 = instruction_io_deq_bits_opcode == 4'h2 ? 4'h0 : _GEN_486; // @[Decoder.scala 373:59]
  wire  _GEN_557 = instruction_io_deq_bits_opcode == 4'h2 ? 1'h0 : _GEN_487; // @[Decoder.scala 373:59]
  wire  _GEN_558 = instruction_io_deq_bits_opcode == 4'h2 ? 1'h0 : _GEN_488; // @[Decoder.scala 373:59]
  wire  _GEN_559 = instruction_io_deq_bits_opcode == 4'h2 ? 1'h0 : _GEN_489; // @[Decoder.scala 373:59]
  wire [11:0] _GEN_560 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_417 : _GEN_490; // @[Decoder.scala 373:59]
  wire [11:0] _GEN_561 = instruction_io_deq_bits_opcode == 4'h2 ? 12'h0 : _GEN_491; // @[Decoder.scala 373:59]
  wire  _GEN_562 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_407 : _GEN_492; // @[Decoder.scala 373:59]
  wire  _GEN_563 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_420 : _GEN_493; // @[Decoder.scala 373:59]
  wire  _GEN_564 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_421 : _GEN_494; // @[Decoder.scala 373:59]
  wire [11:0] _GEN_565 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_422 : 12'h0; // @[Decoder.scala 373:59]
  wire [2:0] _GEN_566 = instruction_io_deq_bits_opcode == 4'h2 ? _GEN_423 : 3'h0; // @[Decoder.scala 373:59]
  wire  _GEN_568 = instruction_io_deq_bits_opcode == 4'h2 ? 1'h0 : _GEN_483; // @[Decoder.scala 373:59 MultiEnqueue.scala 40:17]
  wire  _GEN_569 = instruction_io_deq_bits_opcode == 4'h2 ? 1'h0 : _GEN_484; // @[Decoder.scala 373:59 MultiEnqueue.scala 42:18]
  wire [43:0] _GEN_570 = instruction_io_deq_bits_opcode == 4'h2 ? {{12'd0}, dram0AddressOffset} : _GEN_499; // @[Decoder.scala 126:35 373:59]
  wire [27:0] _GEN_571 = instruction_io_deq_bits_opcode == 4'h2 ? {{24'd0}, dram0CacheBehaviour} : _GEN_500; // @[Decoder.scala 129:36 373:59]
  wire [43:0] _GEN_572 = instruction_io_deq_bits_opcode == 4'h2 ? {{12'd0}, dram1AddressOffset} : _GEN_501; // @[Decoder.scala 130:35 373:59]
  wire [27:0] _GEN_573 = instruction_io_deq_bits_opcode == 4'h2 ? {{24'd0}, dram1CacheBehaviour} : _GEN_502; // @[Decoder.scala 133:36 373:59]
  wire [27:0] _GEN_574 = instruction_io_deq_bits_opcode == 4'h2 ? {{12'd0}, timeout} : _GEN_503; // @[Decoder.scala 373:59 96:24]
  wire  _GEN_580 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_56 : _GEN_568; // @[Decoder.scala 333:62]
  wire  _GEN_581 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_57 : _GEN_569; // @[Decoder.scala 333:62]
  wire  _GEN_582 = instruction_io_deq_bits_opcode == 4'h3 & _GEN_58; // @[Decoder.scala 333:62 670:16]
  wire  _GEN_584 = instruction_io_deq_bits_opcode == 4'h3 & flags_accumulate; // @[Decoder.scala 333:62 669:15]
  wire [13:0] _GEN_585 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_61 : 14'h0; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_586 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_62 : _GEN_539; // @[Decoder.scala 333:62]
  wire  _GEN_587 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_63 : _GEN_509; // @[Decoder.scala 333:62]
  wire  _GEN_588 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_64 : _GEN_510; // @[Decoder.scala 333:62]
  wire  _GEN_589 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_65 : _GEN_546; // @[Decoder.scala 333:62]
  wire [3:0] _GEN_590 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_66 : _GEN_547; // @[Decoder.scala 333:62]
  wire [13:0] _GEN_591 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_67 : _GEN_548; // @[Decoder.scala 333:62]
  wire  _GEN_592 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_68 : _GEN_514; // @[Decoder.scala 333:62]
  wire  _GEN_593 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_69 : _GEN_521; // @[Decoder.scala 333:62]
  wire  _GEN_594 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_70 : _GEN_549; // @[Decoder.scala 333:62]
  wire  _GEN_595 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_550; // @[Decoder.scala 333:62]
  wire [13:0] _GEN_596 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_72 : _GEN_551; // @[Decoder.scala 333:62]
  wire [2:0] _GEN_598 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_74 : _GEN_553; // @[Decoder.scala 333:62]
  wire  _GEN_599 = instruction_io_deq_bits_opcode == 4'h3 & _GEN_75; // @[Decoder.scala 333:62]
  wire  _GEN_600 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_76 : _GEN_528; // @[Decoder.scala 333:62]
  wire  _GEN_601 = instruction_io_deq_bits_opcode == 4'h3 ? _GEN_77 : _GEN_529; // @[Decoder.scala 333:62]
  wire  _GEN_602 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_387; // @[Decoder.scala 333:62]
  wire [13:0] _GEN_603 = instruction_io_deq_bits_opcode == 4'h3 ? req_1_address : args_memAddress; // @[Decoder.scala 333:62]
  wire [13:0] _GEN_604 = instruction_io_deq_bits_opcode == 4'h3 ? instruction_io_deq_ready_w_7_size : _GEN_389; // @[Decoder.scala 333:62]
  wire [2:0] _GEN_605 = instruction_io_deq_bits_opcode == 4'h3 ? args_1_stride : args_memStride; // @[Decoder.scala 333:62]
  wire  _GEN_607 = instruction_io_deq_bits_opcode == 4'h3 ? instruction_io_deq_ready_w_10_lock : _GEN_392; // @[Decoder.scala 333:62]
  wire  _GEN_609 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_394; // @[Decoder.scala 333:62]
  wire  _GEN_611 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_511; // @[Decoder.scala 333:62 670:16]
  wire [1:0] _GEN_612 = instruction_io_deq_bits_opcode == 4'h3 ? 2'h0 : _GEN_512; // @[Decoder.scala 333:62 669:15]
  wire [13:0] _GEN_613 = instruction_io_deq_bits_opcode == 4'h3 ? 14'h0 : _GEN_513; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_614 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_515; // @[Decoder.scala 333:62 670:16]
  wire  _GEN_615 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_516; // @[Decoder.scala 333:62 669:15]
  wire [13:0] _GEN_616 = instruction_io_deq_bits_opcode == 4'h3 ? 14'h0 : _GEN_517; // @[Decoder.scala 333:62 669:15]
  wire [2:0] _GEN_618 = instruction_io_deq_bits_opcode == 4'h3 ? 3'h0 : _GEN_519; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_620 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_522; // @[Decoder.scala 333:62 670:16]
  wire  _GEN_621 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_523; // @[Decoder.scala 333:62 669:15]
  wire [20:0] _GEN_622 = instruction_io_deq_bits_opcode == 4'h3 ? 21'h0 : _GEN_524; // @[Decoder.scala 333:62 669:15]
  wire [20:0] _GEN_623 = instruction_io_deq_bits_opcode == 4'h3 ? 21'h0 : _GEN_525; // @[Decoder.scala 333:62 669:15]
  wire [2:0] _GEN_624 = instruction_io_deq_bits_opcode == 4'h3 ? 3'h0 : _GEN_526; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_626 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_540; // @[Decoder.scala 333:62 670:16]
  wire  _GEN_627 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_541; // @[Decoder.scala 333:62 669:15]
  wire [20:0] _GEN_628 = instruction_io_deq_bits_opcode == 4'h3 ? 21'h0 : _GEN_542; // @[Decoder.scala 333:62 669:15]
  wire [20:0] _GEN_629 = instruction_io_deq_bits_opcode == 4'h3 ? 21'h0 : _GEN_543; // @[Decoder.scala 333:62 669:15]
  wire [2:0] _GEN_630 = instruction_io_deq_bits_opcode == 4'h3 ? 3'h0 : _GEN_544; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_632 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_555; // @[Decoder.scala 333:62 670:16]
  wire [3:0] _GEN_633 = instruction_io_deq_bits_opcode == 4'h3 ? 4'h0 : _GEN_556; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_634 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_557; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_635 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_558; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_636 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_559; // @[Decoder.scala 333:62 669:15]
  wire [11:0] _GEN_637 = instruction_io_deq_bits_opcode == 4'h3 ? 12'h0 : _GEN_560; // @[Decoder.scala 333:62 669:15]
  wire [11:0] _GEN_638 = instruction_io_deq_bits_opcode == 4'h3 ? 12'h0 : _GEN_561; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_639 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_562; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_640 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_563; // @[Decoder.scala 333:62 669:15]
  wire  _GEN_641 = instruction_io_deq_bits_opcode == 4'h3 ? 1'h0 : _GEN_564; // @[Decoder.scala 333:62 669:15]
  wire [11:0] _GEN_642 = instruction_io_deq_bits_opcode == 4'h3 ? 12'h0 : _GEN_565; // @[Decoder.scala 333:62 669:15]
  wire [2:0] _GEN_643 = instruction_io_deq_bits_opcode == 4'h3 ? 3'h0 : _GEN_566; // @[Decoder.scala 333:62 669:15]
  wire [43:0] _GEN_645 = instruction_io_deq_bits_opcode == 4'h3 ? {{12'd0}, dram0AddressOffset} : _GEN_570; // @[Decoder.scala 126:35 333:62]
  wire [27:0] _GEN_646 = instruction_io_deq_bits_opcode == 4'h3 ? {{24'd0}, dram0CacheBehaviour} : _GEN_571; // @[Decoder.scala 129:36 333:62]
  wire [43:0] _GEN_647 = instruction_io_deq_bits_opcode == 4'h3 ? {{12'd0}, dram1AddressOffset} : _GEN_572; // @[Decoder.scala 130:35 333:62]
  wire [27:0] _GEN_648 = instruction_io_deq_bits_opcode == 4'h3 ? {{24'd0}, dram1CacheBehaviour} : _GEN_573; // @[Decoder.scala 133:36 333:62]
  wire [27:0] _GEN_649 = instruction_io_deq_bits_opcode == 4'h3 ? {{12'd0}, timeout} : _GEN_574; // @[Decoder.scala 333:62 96:24]
  wire [43:0] _GEN_730 = instruction_io_deq_bits_opcode == 4'h1 ? {{12'd0}, dram0AddressOffset} : _GEN_645; // @[Decoder.scala 126:35 282:51]
  wire [27:0] _GEN_731 = instruction_io_deq_bits_opcode == 4'h1 ? {{24'd0}, dram0CacheBehaviour} : _GEN_646; // @[Decoder.scala 129:36 282:51]
  wire [43:0] _GEN_732 = instruction_io_deq_bits_opcode == 4'h1 ? {{12'd0}, dram1AddressOffset} : _GEN_647; // @[Decoder.scala 130:35 282:51]
  wire [27:0] _GEN_733 = instruction_io_deq_bits_opcode == 4'h1 ? {{24'd0}, dram1CacheBehaviour} : _GEN_648; // @[Decoder.scala 133:36 282:51]
  wire [27:0] _GEN_734 = instruction_io_deq_bits_opcode == 4'h1 ? {{12'd0}, timeout} : _GEN_649; // @[Decoder.scala 282:51 96:24]
  wire [27:0] _GEN_86 = reset ? 28'h64 : _GEN_734; // @[Decoder.scala 96:{24,24}]
  wire [43:0] _GEN_123 = reset ? 44'h0 : _GEN_730; // @[Decoder.scala 126:{35,35}]
  wire [27:0] _GEN_161 = reset ? 28'h0 : _GEN_731; // @[Decoder.scala 129:{36,36}]
  wire [43:0] _GEN_199 = reset ? 44'h0 : _GEN_732; // @[Decoder.scala 130:{35,35}]
  wire [27:0] _GEN_230 = reset ? 28'h0 : _GEN_733; // @[Decoder.scala 133:{36,36}]
  Queue instruction ( // @[Decoupled.scala 361:21]
    .clock(instruction_clock),
    .reset(instruction_reset),
    .io_enq_ready(instruction_io_enq_ready),
    .io_enq_valid(instruction_io_enq_valid),
    .io_enq_bits_opcode(instruction_io_enq_bits_opcode),
    .io_enq_bits_flags(instruction_io_enq_bits_flags),
    .io_enq_bits_arguments(instruction_io_enq_bits_arguments),
    .io_deq_ready(instruction_io_deq_ready),
    .io_deq_valid(instruction_io_deq_valid),
    .io_deq_bits_opcode(instruction_io_deq_bits_opcode),
    .io_deq_bits_flags(instruction_io_deq_bits_flags),
    .io_deq_bits_arguments(instruction_io_deq_bits_arguments)
  );
  StrideHandler dram0Handler ( // @[Decoder.scala 144:28]
    .clock(dram0Handler_clock),
    .reset(dram0Handler_reset),
    .io_in_ready(dram0Handler_io_in_ready),
    .io_in_valid(dram0Handler_io_in_valid),
    .io_in_bits_write(dram0Handler_io_in_bits_write),
    .io_in_bits_address(dram0Handler_io_in_bits_address),
    .io_in_bits_size(dram0Handler_io_in_bits_size),
    .io_in_bits_stride(dram0Handler_io_in_bits_stride),
    .io_in_bits_reverse(dram0Handler_io_in_bits_reverse),
    .io_out_ready(dram0Handler_io_out_ready),
    .io_out_valid(dram0Handler_io_out_valid),
    .io_out_bits_write(dram0Handler_io_out_bits_write),
    .io_out_bits_address(dram0Handler_io_out_bits_address),
    .io_out_bits_size(dram0Handler_io_out_bits_size)
  );
  StrideHandler dram1Handler ( // @[Decoder.scala 153:28]
    .clock(dram1Handler_clock),
    .reset(dram1Handler_reset),
    .io_in_ready(dram1Handler_io_in_ready),
    .io_in_valid(dram1Handler_io_in_valid),
    .io_in_bits_write(dram1Handler_io_in_bits_write),
    .io_in_bits_address(dram1Handler_io_in_bits_address),
    .io_in_bits_size(dram1Handler_io_in_bits_size),
    .io_in_bits_stride(dram1Handler_io_in_bits_stride),
    .io_in_bits_reverse(dram1Handler_io_in_bits_reverse),
    .io_out_ready(dram1Handler_io_out_ready),
    .io_out_valid(dram1Handler_io_out_valid),
    .io_out_bits_write(dram1Handler_io_out_bits_write),
    .io_out_bits_address(dram1Handler_io_out_bits_address),
    .io_out_bits_size(dram1Handler_io_out_bits_size)
  );
  Queue_2 dram0 ( // @[Mem.scala 22:19]
    .clock(dram0_clock),
    .reset(dram0_reset),
    .io_enq_ready(dram0_io_enq_ready),
    .io_enq_valid(dram0_io_enq_valid),
    .io_enq_bits_write(dram0_io_enq_bits_write),
    .io_enq_bits_address(dram0_io_enq_bits_address),
    .io_enq_bits_size(dram0_io_enq_bits_size),
    .io_enq_bits_stride(dram0_io_enq_bits_stride),
    .io_deq_ready(dram0_io_deq_ready),
    .io_deq_valid(dram0_io_deq_valid),
    .io_deq_bits_write(dram0_io_deq_bits_write),
    .io_deq_bits_address(dram0_io_deq_bits_address),
    .io_deq_bits_size(dram0_io_deq_bits_size),
    .io_deq_bits_stride(dram0_io_deq_bits_stride),
    .io_deq_bits_reverse(dram0_io_deq_bits_reverse)
  );
  Queue_2 dram1 ( // @[Mem.scala 22:19]
    .clock(dram1_clock),
    .reset(dram1_reset),
    .io_enq_ready(dram1_io_enq_ready),
    .io_enq_valid(dram1_io_enq_valid),
    .io_enq_bits_write(dram1_io_enq_bits_write),
    .io_enq_bits_address(dram1_io_enq_bits_address),
    .io_enq_bits_size(dram1_io_enq_bits_size),
    .io_enq_bits_stride(dram1_io_enq_bits_stride),
    .io_deq_ready(dram1_io_deq_ready),
    .io_deq_valid(dram1_io_deq_valid),
    .io_deq_bits_write(dram1_io_deq_bits_write),
    .io_deq_bits_address(dram1_io_deq_bits_address),
    .io_deq_bits_size(dram1_io_deq_bits_size),
    .io_deq_bits_stride(dram1_io_deq_bits_stride),
    .io_deq_bits_reverse(dram1_io_deq_bits_reverse)
  );
  SizeAndStrideHandler_2 memPortAHandler ( // @[Decoder.scala 168:31]
    .clock(memPortAHandler_clock),
    .reset(memPortAHandler_reset),
    .io_in_ready(memPortAHandler_io_in_ready),
    .io_in_valid(memPortAHandler_io_in_valid),
    .io_in_bits_write(memPortAHandler_io_in_bits_write),
    .io_in_bits_address(memPortAHandler_io_in_bits_address),
    .io_in_bits_size(memPortAHandler_io_in_bits_size),
    .io_in_bits_stride(memPortAHandler_io_in_bits_stride),
    .io_in_bits_reverse(memPortAHandler_io_in_bits_reverse),
    .io_out_ready(memPortAHandler_io_out_ready),
    .io_out_valid(memPortAHandler_io_out_valid),
    .io_out_bits_write(memPortAHandler_io_out_bits_write),
    .io_out_bits_address(memPortAHandler_io_out_bits_address)
  );
  SizeAndStrideHandler_2 memPortBHandler ( // @[Decoder.scala 177:31]
    .clock(memPortBHandler_clock),
    .reset(memPortBHandler_reset),
    .io_in_ready(memPortBHandler_io_in_ready),
    .io_in_valid(memPortBHandler_io_in_valid),
    .io_in_bits_write(memPortBHandler_io_in_bits_write),
    .io_in_bits_address(memPortBHandler_io_in_bits_address),
    .io_in_bits_size(memPortBHandler_io_in_bits_size),
    .io_in_bits_stride(memPortBHandler_io_in_bits_stride),
    .io_in_bits_reverse(memPortBHandler_io_in_bits_reverse),
    .io_out_ready(memPortBHandler_io_out_ready),
    .io_out_valid(memPortBHandler_io_out_valid),
    .io_out_bits_write(memPortBHandler_io_out_bits_write),
    .io_out_bits_address(memPortBHandler_io_out_bits_address)
  );
  LockPool lockPool ( // @[Decoder.scala 193:24]
    .clock(lockPool_clock),
    .reset(lockPool_reset),
    .io_actor_0_in_ready(lockPool_io_actor_0_in_ready),
    .io_actor_0_in_valid(lockPool_io_actor_0_in_valid),
    .io_actor_0_in_bits_write(lockPool_io_actor_0_in_bits_write),
    .io_actor_0_in_bits_address(lockPool_io_actor_0_in_bits_address),
    .io_actor_0_in_bits_size(lockPool_io_actor_0_in_bits_size),
    .io_actor_0_in_bits_stride(lockPool_io_actor_0_in_bits_stride),
    .io_actor_0_in_bits_reverse(lockPool_io_actor_0_in_bits_reverse),
    .io_actor_0_out_ready(lockPool_io_actor_0_out_ready),
    .io_actor_0_out_valid(lockPool_io_actor_0_out_valid),
    .io_actor_0_out_bits_write(lockPool_io_actor_0_out_bits_write),
    .io_actor_0_out_bits_address(lockPool_io_actor_0_out_bits_address),
    .io_actor_0_out_bits_size(lockPool_io_actor_0_out_bits_size),
    .io_actor_0_out_bits_stride(lockPool_io_actor_0_out_bits_stride),
    .io_actor_0_out_bits_reverse(lockPool_io_actor_0_out_bits_reverse),
    .io_actor_1_in_ready(lockPool_io_actor_1_in_ready),
    .io_actor_1_in_valid(lockPool_io_actor_1_in_valid),
    .io_actor_1_in_bits_write(lockPool_io_actor_1_in_bits_write),
    .io_actor_1_in_bits_address(lockPool_io_actor_1_in_bits_address),
    .io_actor_1_in_bits_size(lockPool_io_actor_1_in_bits_size),
    .io_actor_1_in_bits_stride(lockPool_io_actor_1_in_bits_stride),
    .io_actor_1_out_ready(lockPool_io_actor_1_out_ready),
    .io_actor_1_out_valid(lockPool_io_actor_1_out_valid),
    .io_actor_1_out_bits_write(lockPool_io_actor_1_out_bits_write),
    .io_actor_1_out_bits_address(lockPool_io_actor_1_out_bits_address),
    .io_actor_1_out_bits_size(lockPool_io_actor_1_out_bits_size),
    .io_actor_1_out_bits_stride(lockPool_io_actor_1_out_bits_stride),
    .io_actor_1_out_bits_reverse(lockPool_io_actor_1_out_bits_reverse),
    .io_lock_ready(lockPool_io_lock_ready),
    .io_lock_valid(lockPool_io_lock_valid),
    .io_lock_bits_cond_write(lockPool_io_lock_bits_cond_write),
    .io_lock_bits_cond_address(lockPool_io_lock_bits_cond_address),
    .io_lock_bits_cond_size(lockPool_io_lock_bits_cond_size),
    .io_lock_bits_cond_stride(lockPool_io_lock_bits_cond_stride),
    .io_lock_bits_cond_reverse(lockPool_io_lock_bits_cond_reverse),
    .io_lock_bits_lock(lockPool_io_lock_bits_lock),
    .io_lock_bits_by(lockPool_io_lock_bits_by)
  );
  SizeAndStrideHandler_4 accHandler ( // @[Decoder.scala 207:26]
    .clock(accHandler_clock),
    .reset(accHandler_reset),
    .io_in_ready(accHandler_io_in_ready),
    .io_in_valid(accHandler_io_in_valid),
    .io_in_bits_instruction_op(accHandler_io_in_bits_instruction_op),
    .io_in_bits_instruction_sourceLeft(accHandler_io_in_bits_instruction_sourceLeft),
    .io_in_bits_instruction_sourceRight(accHandler_io_in_bits_instruction_sourceRight),
    .io_in_bits_instruction_dest(accHandler_io_in_bits_instruction_dest),
    .io_in_bits_address(accHandler_io_in_bits_address),
    .io_in_bits_altAddress(accHandler_io_in_bits_altAddress),
    .io_in_bits_read(accHandler_io_in_bits_read),
    .io_in_bits_write(accHandler_io_in_bits_write),
    .io_in_bits_accumulate(accHandler_io_in_bits_accumulate),
    .io_in_bits_size(accHandler_io_in_bits_size),
    .io_in_bits_stride(accHandler_io_in_bits_stride),
    .io_in_bits_reverse(accHandler_io_in_bits_reverse),
    .io_out_ready(accHandler_io_out_ready),
    .io_out_valid(accHandler_io_out_valid),
    .io_out_bits_instruction_op(accHandler_io_out_bits_instruction_op),
    .io_out_bits_instruction_sourceLeft(accHandler_io_out_bits_instruction_sourceLeft),
    .io_out_bits_instruction_sourceRight(accHandler_io_out_bits_instruction_sourceRight),
    .io_out_bits_instruction_dest(accHandler_io_out_bits_instruction_dest),
    .io_out_bits_address(accHandler_io_out_bits_address),
    .io_out_bits_altAddress(accHandler_io_out_bits_altAddress),
    .io_out_bits_read(accHandler_io_out_bits_read),
    .io_out_bits_write(accHandler_io_out_bits_write),
    .io_out_bits_accumulate(accHandler_io_out_bits_accumulate)
  );
  Queue_4 acc ( // @[Mem.scala 22:19]
    .clock(acc_clock),
    .reset(acc_reset),
    .io_enq_ready(acc_io_enq_ready),
    .io_enq_valid(acc_io_enq_valid),
    .io_enq_bits_instruction_op(acc_io_enq_bits_instruction_op),
    .io_enq_bits_instruction_sourceLeft(acc_io_enq_bits_instruction_sourceLeft),
    .io_enq_bits_instruction_sourceRight(acc_io_enq_bits_instruction_sourceRight),
    .io_enq_bits_instruction_dest(acc_io_enq_bits_instruction_dest),
    .io_enq_bits_address(acc_io_enq_bits_address),
    .io_enq_bits_altAddress(acc_io_enq_bits_altAddress),
    .io_enq_bits_read(acc_io_enq_bits_read),
    .io_enq_bits_write(acc_io_enq_bits_write),
    .io_enq_bits_accumulate(acc_io_enq_bits_accumulate),
    .io_enq_bits_size(acc_io_enq_bits_size),
    .io_enq_bits_stride(acc_io_enq_bits_stride),
    .io_deq_ready(acc_io_deq_ready),
    .io_deq_valid(acc_io_deq_valid),
    .io_deq_bits_instruction_op(acc_io_deq_bits_instruction_op),
    .io_deq_bits_instruction_sourceLeft(acc_io_deq_bits_instruction_sourceLeft),
    .io_deq_bits_instruction_sourceRight(acc_io_deq_bits_instruction_sourceRight),
    .io_deq_bits_instruction_dest(acc_io_deq_bits_instruction_dest),
    .io_deq_bits_address(acc_io_deq_bits_address),
    .io_deq_bits_altAddress(acc_io_deq_bits_altAddress),
    .io_deq_bits_read(acc_io_deq_bits_read),
    .io_deq_bits_write(acc_io_deq_bits_write),
    .io_deq_bits_accumulate(acc_io_deq_bits_accumulate),
    .io_deq_bits_size(acc_io_deq_bits_size),
    .io_deq_bits_stride(acc_io_deq_bits_stride),
    .io_deq_bits_reverse(acc_io_deq_bits_reverse)
  );
  SizeHandler arrayHandler ( // @[Decoder.scala 230:28]
    .clock(arrayHandler_clock),
    .reset(arrayHandler_reset),
    .io_in_ready(arrayHandler_io_in_ready),
    .io_in_valid(arrayHandler_io_in_valid),
    .io_in_bits_load(arrayHandler_io_in_bits_load),
    .io_in_bits_zeroes(arrayHandler_io_in_bits_zeroes),
    .io_in_bits_size(arrayHandler_io_in_bits_size),
    .io_out_ready(arrayHandler_io_out_ready),
    .io_out_valid(arrayHandler_io_out_valid),
    .io_out_bits_load(arrayHandler_io_out_bits_load),
    .io_out_bits_zeroes(arrayHandler_io_out_bits_zeroes)
  );
  Queue_5 array ( // @[Mem.scala 22:19]
    .clock(array_clock),
    .reset(array_reset),
    .io_enq_ready(array_io_enq_ready),
    .io_enq_valid(array_io_enq_valid),
    .io_enq_bits_load(array_io_enq_bits_load),
    .io_enq_bits_zeroes(array_io_enq_bits_zeroes),
    .io_enq_bits_size(array_io_enq_bits_size),
    .io_deq_ready(array_io_deq_ready),
    .io_deq_valid(array_io_deq_valid),
    .io_deq_bits_load(array_io_deq_bits_load),
    .io_deq_bits_zeroes(array_io_deq_bits_zeroes),
    .io_deq_bits_size(array_io_deq_bits_size)
  );
  Queue_6 dataflow ( // @[Mem.scala 22:19]
    .clock(dataflow_clock),
    .reset(dataflow_reset),
    .io_enq_ready(dataflow_io_enq_ready),
    .io_enq_valid(dataflow_io_enq_valid),
    .io_enq_bits_kind(dataflow_io_enq_bits_kind),
    .io_enq_bits_size(dataflow_io_enq_bits_size),
    .io_deq_ready(dataflow_io_deq_ready),
    .io_deq_valid(dataflow_io_deq_valid),
    .io_deq_bits_kind(dataflow_io_deq_bits_kind),
    .io_deq_bits_size(dataflow_io_deq_bits_size)
  );
  SizeHandler_1 hostDataflowHandler ( // @[Decoder.scala 250:35]
    .clock(hostDataflowHandler_clock),
    .reset(hostDataflowHandler_reset),
    .io_in_ready(hostDataflowHandler_io_in_ready),
    .io_in_valid(hostDataflowHandler_io_in_valid),
    .io_in_bits_kind(hostDataflowHandler_io_in_bits_kind),
    .io_in_bits_size(hostDataflowHandler_io_in_bits_size),
    .io_out_ready(hostDataflowHandler_io_out_ready),
    .io_out_valid(hostDataflowHandler_io_out_valid),
    .io_out_bits_kind(hostDataflowHandler_io_out_bits_kind)
  );
  Queue_7 hostDataflow ( // @[Mem.scala 22:19]
    .clock(hostDataflow_clock),
    .reset(hostDataflow_reset),
    .io_enq_ready(hostDataflow_io_enq_ready),
    .io_enq_valid(hostDataflow_io_enq_valid),
    .io_enq_bits_kind(hostDataflow_io_enq_bits_kind),
    .io_enq_bits_size(hostDataflow_io_enq_bits_size),
    .io_deq_ready(hostDataflow_io_deq_ready),
    .io_deq_valid(hostDataflow_io_deq_valid),
    .io_deq_bits_kind(hostDataflow_io_deq_bits_kind),
    .io_deq_bits_size(hostDataflow_io_deq_bits_size)
  );
  MultiEnqueue enqueuer1 ( // @[MultiEnqueue.scala 182:43]
    .clock(enqueuer1_clock),
    .reset(enqueuer1_reset),
    .io_in_ready(enqueuer1_io_in_ready),
    .io_in_valid(enqueuer1_io_in_valid),
    .io_out_0_ready(enqueuer1_io_out_0_ready),
    .io_out_0_valid(enqueuer1_io_out_0_valid)
  );
  MultiEnqueue_1 enqueuer2 ( // @[MultiEnqueue.scala 182:43]
    .clock(enqueuer2_clock),
    .reset(enqueuer2_reset),
    .io_in_ready(enqueuer2_io_in_ready),
    .io_in_valid(enqueuer2_io_in_valid),
    .io_out_0_ready(enqueuer2_io_out_0_ready),
    .io_out_0_valid(enqueuer2_io_out_0_valid),
    .io_out_1_ready(enqueuer2_io_out_1_ready),
    .io_out_1_valid(enqueuer2_io_out_1_valid)
  );
  MultiEnqueue_2 enqueuer3 ( // @[MultiEnqueue.scala 182:43]
    .clock(enqueuer3_clock),
    .reset(enqueuer3_reset),
    .io_in_ready(enqueuer3_io_in_ready),
    .io_in_valid(enqueuer3_io_in_valid),
    .io_out_0_ready(enqueuer3_io_out_0_ready),
    .io_out_0_valid(enqueuer3_io_out_0_valid),
    .io_out_1_ready(enqueuer3_io_out_1_ready),
    .io_out_1_valid(enqueuer3_io_out_1_valid),
    .io_out_2_ready(enqueuer3_io_out_2_ready),
    .io_out_2_valid(enqueuer3_io_out_2_valid)
  );
  MultiEnqueue_3 enqueuer4 ( // @[MultiEnqueue.scala 182:43]
    .clock(enqueuer4_clock),
    .reset(enqueuer4_reset),
    .io_in_ready(enqueuer4_io_in_ready),
    .io_in_valid(enqueuer4_io_in_valid),
    .io_out_0_ready(enqueuer4_io_out_0_ready),
    .io_out_0_valid(enqueuer4_io_out_0_valid),
    .io_out_1_ready(enqueuer4_io_out_1_ready),
    .io_out_1_valid(enqueuer4_io_out_1_valid),
    .io_out_2_ready(enqueuer4_io_out_2_ready),
    .io_out_2_valid(enqueuer4_io_out_2_valid),
    .io_out_3_ready(enqueuer4_io_out_3_ready),
    .io_out_3_valid(enqueuer4_io_out_3_valid)
  );
  MultiEnqueue_4 enqueuer5 ( // @[MultiEnqueue.scala 182:43]
    .clock(enqueuer5_clock),
    .reset(enqueuer5_reset),
    .io_in_ready(enqueuer5_io_in_ready),
    .io_in_valid(enqueuer5_io_in_valid),
    .io_out_0_ready(enqueuer5_io_out_0_ready),
    .io_out_0_valid(enqueuer5_io_out_0_valid),
    .io_out_1_ready(enqueuer5_io_out_1_ready),
    .io_out_1_valid(enqueuer5_io_out_1_valid),
    .io_out_2_ready(enqueuer5_io_out_2_ready),
    .io_out_2_valid(enqueuer5_io_out_2_valid),
    .io_out_3_ready(enqueuer5_io_out_3_ready),
    .io_out_3_valid(enqueuer5_io_out_3_valid),
    .io_out_4_ready(enqueuer5_io_out_4_ready),
    .io_out_4_valid(enqueuer5_io_out_4_valid)
  );
  assign io_instruction_ready = instruction_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_memPortA_valid = memPortAHandler_io_out_valid; // @[Decoder.scala 186:15]
  assign io_memPortA_bits_write = memPortAHandler_io_out_bits_write; // @[Decoder.scala 186:15]
  assign io_memPortA_bits_address = memPortAHandler_io_out_bits_address; // @[Decoder.scala 186:15]
  assign io_memPortB_valid = memPortBHandler_io_out_valid; // @[Decoder.scala 187:15]
  assign io_memPortB_bits_write = memPortBHandler_io_out_bits_write; // @[Decoder.scala 187:15]
  assign io_memPortB_bits_address = memPortBHandler_io_out_bits_address; // @[Decoder.scala 187:15]
  assign io_dram0_valid = dram0Handler_io_out_valid; // @[Decoder.scala 162:12]
  assign io_dram0_bits_write = dram0Handler_io_out_bits_write; // @[Decoder.scala 162:12]
  assign io_dram0_bits_address = dram0Handler_io_out_bits_address; // @[Decoder.scala 162:12]
  assign io_dram0_bits_size = dram0Handler_io_out_bits_size; // @[Decoder.scala 162:12]
  assign io_dram1_valid = dram1Handler_io_out_valid; // @[Decoder.scala 163:12]
  assign io_dram1_bits_write = dram1Handler_io_out_bits_write; // @[Decoder.scala 163:12]
  assign io_dram1_bits_address = dram1Handler_io_out_bits_address; // @[Decoder.scala 163:12]
  assign io_dram1_bits_size = dram1Handler_io_out_bits_size; // @[Decoder.scala 163:12]
  assign io_dataflow_valid = dataflow_io_deq_valid; // @[Mem.scala 23:7]
  assign io_dataflow_bits_kind = dataflow_io_deq_bits_kind; // @[Mem.scala 23:7]
  assign io_dataflow_bits_size = dataflow_io_deq_bits_size; // @[Mem.scala 23:7]
  assign io_hostDataflow_valid = hostDataflowHandler_io_out_valid; // @[Decoder.scala 257:19]
  assign io_hostDataflow_bits_kind = hostDataflowHandler_io_out_bits_kind; // @[Decoder.scala 257:19]
  assign io_acc_valid = accHandler_io_out_valid; // @[Decoder.scala 218:16]
  assign io_acc_bits_instruction_op = accHandler_io_out_bits_instruction_op; // @[AccumulatorWithALUArrayControl.scala 96:17 102:19]
  assign io_acc_bits_instruction_sourceLeft = accHandler_io_out_bits_instruction_sourceLeft; // @[AccumulatorWithALUArrayControl.scala 96:17 102:19]
  assign io_acc_bits_instruction_sourceRight = accHandler_io_out_bits_instruction_sourceRight; // @[AccumulatorWithALUArrayControl.scala 96:17 102:19]
  assign io_acc_bits_instruction_dest = accHandler_io_out_bits_instruction_dest; // @[AccumulatorWithALUArrayControl.scala 96:17 102:19]
  assign io_acc_bits_readAddress = io_acc_bits_isMemControl ? _GEN_5 : accHandler_io_out_bits_address; // @[AccumulatorWithALUArrayControl.scala 106:24 120:21]
  assign io_acc_bits_writeAddress = io_acc_bits_isMemControl ? _GEN_6 : accHandler_io_out_bits_altAddress; // @[AccumulatorWithALUArrayControl.scala 106:24 121:22]
  assign io_acc_bits_accumulate = accHandler_io_out_bits_accumulate; // @[AccumulatorWithALUArrayControl.scala 96:17 105:18]
  assign io_acc_bits_write = accHandler_io_out_bits_write; // @[AccumulatorWithALUArrayControl.scala 104:13 96:17]
  assign io_acc_bits_read = accHandler_io_out_bits_read; // @[AccumulatorWithALUArrayControl.scala 103:12 96:17]
  assign io_array_valid = arrayHandler_io_out_valid; // @[Decoder.scala 239:12]
  assign io_array_bits_load = arrayHandler_io_out_bits_load; // @[Decoder.scala 239:12]
  assign io_array_bits_zeroes = arrayHandler_io_out_bits_zeroes; // @[Decoder.scala 239:12]
  assign io_config_dram0AddressOffset = dram0AddressOffset; // @[Decoder.scala 135:32]
  assign io_config_dram0CacheBehaviour = dram0CacheBehaviour; // @[Decoder.scala 136:33]
  assign io_config_dram1AddressOffset = dram1AddressOffset; // @[Decoder.scala 137:32]
  assign io_config_dram1CacheBehaviour = dram1CacheBehaviour; // @[Decoder.scala 138:33]
  assign io_timeout = timer == timeout; // @[Decoder.scala 105:23]
  assign io_error = 1'h0; // @[Decoder.scala 646:14]
  assign io_tracepoint = programCounter == tracepoint; // @[Decoder.scala 113:35]
  assign io_programCounter = programCounter; // @[Decoder.scala 114:21]
  assign instruction_clock = clock;
  assign instruction_reset = reset;
  assign instruction_io_enq_valid = io_instruction_valid; // @[Decoupled.scala 363:22]
  assign instruction_io_enq_bits_opcode = io_instruction_bits_opcode; // @[Decoupled.scala 364:21]
  assign instruction_io_enq_bits_flags = io_instruction_bits_flags; // @[Decoupled.scala 364:21]
  assign instruction_io_enq_bits_arguments = io_instruction_bits_arguments; // @[Decoupled.scala 364:21]
  assign instruction_io_deq_ready = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_33 : _GEN_586; // @[Decoder.scala 282:51]
  assign dram0Handler_clock = clock;
  assign dram0Handler_reset = reset;
  assign dram0Handler_io_in_valid = dram0_io_deq_valid; // @[Mem.scala 23:7]
  assign dram0Handler_io_in_bits_write = dram0_io_deq_bits_write; // @[Mem.scala 23:7]
  assign dram0Handler_io_in_bits_address = dram0_io_deq_bits_address; // @[Mem.scala 23:7]
  assign dram0Handler_io_in_bits_size = dram0_io_deq_bits_size; // @[Mem.scala 23:7]
  assign dram0Handler_io_in_bits_stride = dram0_io_deq_bits_stride; // @[Mem.scala 23:7]
  assign dram0Handler_io_in_bits_reverse = dram0_io_deq_bits_reverse; // @[Mem.scala 23:7]
  assign dram0Handler_io_out_ready = io_dram0_ready; // @[Decoder.scala 162:12]
  assign dram1Handler_clock = clock;
  assign dram1Handler_reset = reset;
  assign dram1Handler_io_in_valid = dram1_io_deq_valid; // @[Mem.scala 23:7]
  assign dram1Handler_io_in_bits_write = dram1_io_deq_bits_write; // @[Mem.scala 23:7]
  assign dram1Handler_io_in_bits_address = dram1_io_deq_bits_address; // @[Mem.scala 23:7]
  assign dram1Handler_io_in_bits_size = dram1_io_deq_bits_size; // @[Mem.scala 23:7]
  assign dram1Handler_io_in_bits_stride = dram1_io_deq_bits_stride; // @[Mem.scala 23:7]
  assign dram1Handler_io_in_bits_reverse = dram1_io_deq_bits_reverse; // @[Mem.scala 23:7]
  assign dram1Handler_io_out_ready = io_dram1_ready; // @[Decoder.scala 163:12]
  assign dram0_clock = clock;
  assign dram0_reset = reset;
  assign dram0_io_enq_valid = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_620; // @[Decoder.scala 282:51 670:16]
  assign dram0_io_enq_bits_write = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_621; // @[Decoder.scala 282:51 669:15]
  assign dram0_io_enq_bits_address = instruction_io_deq_bits_opcode == 4'h1 ? 21'h0 : _GEN_622; // @[Decoder.scala 282:51 669:15]
  assign dram0_io_enq_bits_size = instruction_io_deq_bits_opcode == 4'h1 ? 21'h0 : _GEN_623; // @[Decoder.scala 282:51 669:15]
  assign dram0_io_enq_bits_stride = instruction_io_deq_bits_opcode == 4'h1 ? 3'h0 : _GEN_624; // @[Decoder.scala 282:51 669:15]
  assign dram0_io_deq_ready = dram0Handler_io_in_ready; // @[Mem.scala 23:7]
  assign dram1_clock = clock;
  assign dram1_reset = reset;
  assign dram1_io_enq_valid = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_626; // @[Decoder.scala 282:51 670:16]
  assign dram1_io_enq_bits_write = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_627; // @[Decoder.scala 282:51 669:15]
  assign dram1_io_enq_bits_address = instruction_io_deq_bits_opcode == 4'h1 ? 21'h0 : _GEN_628; // @[Decoder.scala 282:51 669:15]
  assign dram1_io_enq_bits_size = instruction_io_deq_bits_opcode == 4'h1 ? 21'h0 : _GEN_629; // @[Decoder.scala 282:51 669:15]
  assign dram1_io_enq_bits_stride = instruction_io_deq_bits_opcode == 4'h1 ? 3'h0 : _GEN_630; // @[Decoder.scala 282:51 669:15]
  assign dram1_io_deq_ready = dram1Handler_io_in_ready; // @[Mem.scala 23:7]
  assign memPortAHandler_clock = clock;
  assign memPortAHandler_reset = reset;
  assign memPortAHandler_io_in_valid = lockPool_io_actor_0_out_valid; // @[Decoder.scala 196:25]
  assign memPortAHandler_io_in_bits_write = lockPool_io_actor_0_out_bits_write; // @[Decoder.scala 196:25]
  assign memPortAHandler_io_in_bits_address = lockPool_io_actor_0_out_bits_address; // @[Decoder.scala 196:25]
  assign memPortAHandler_io_in_bits_size = lockPool_io_actor_0_out_bits_size; // @[Decoder.scala 196:25]
  assign memPortAHandler_io_in_bits_stride = lockPool_io_actor_0_out_bits_stride; // @[Decoder.scala 196:25]
  assign memPortAHandler_io_in_bits_reverse = lockPool_io_actor_0_out_bits_reverse; // @[Decoder.scala 196:25]
  assign memPortAHandler_io_out_ready = io_memPortA_ready; // @[Decoder.scala 186:15]
  assign memPortBHandler_clock = clock;
  assign memPortBHandler_reset = reset;
  assign memPortBHandler_io_in_valid = lockPool_io_actor_1_out_valid; // @[Decoder.scala 197:25]
  assign memPortBHandler_io_in_bits_write = lockPool_io_actor_1_out_bits_write; // @[Decoder.scala 197:25]
  assign memPortBHandler_io_in_bits_address = lockPool_io_actor_1_out_bits_address; // @[Decoder.scala 197:25]
  assign memPortBHandler_io_in_bits_size = lockPool_io_actor_1_out_bits_size; // @[Decoder.scala 197:25]
  assign memPortBHandler_io_in_bits_stride = lockPool_io_actor_1_out_bits_stride; // @[Decoder.scala 197:25]
  assign memPortBHandler_io_in_bits_reverse = lockPool_io_actor_1_out_bits_reverse; // @[Decoder.scala 197:25]
  assign memPortBHandler_io_out_ready = io_memPortB_ready; // @[Decoder.scala 187:15]
  assign lockPool_clock = clock;
  assign lockPool_reset = reset;
  assign lockPool_io_actor_0_in_valid = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_37 : _GEN_594; // @[Decoder.scala 282:51]
  assign lockPool_io_actor_0_in_bits_write = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_595; // @[Decoder.scala 282:51]
  assign lockPool_io_actor_0_in_bits_address = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_39 : _GEN_596; // @[Decoder.scala 282:51]
  assign lockPool_io_actor_0_in_bits_size = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_40 : _GEN_591; // @[Decoder.scala 282:51]
  assign lockPool_io_actor_0_in_bits_stride = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_41 : _GEN_598; // @[Decoder.scala 282:51]
  assign lockPool_io_actor_0_in_bits_reverse = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_599; // @[Decoder.scala 282:51]
  assign lockPool_io_actor_0_out_ready = memPortAHandler_io_in_ready; // @[Decoder.scala 196:25]
  assign lockPool_io_actor_1_in_valid = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_614; // @[Decoder.scala 282:51 670:16]
  assign lockPool_io_actor_1_in_bits_write = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_615; // @[Decoder.scala 282:51 669:15]
  assign lockPool_io_actor_1_in_bits_address = instruction_io_deq_bits_opcode == 4'h1 ? 14'h0 : _GEN_616; // @[Decoder.scala 282:51 669:15]
  assign lockPool_io_actor_1_in_bits_size = instruction_io_deq_bits_opcode == 4'h1 ? 14'h0 : _GEN_613; // @[Decoder.scala 282:51 669:15]
  assign lockPool_io_actor_1_in_bits_stride = instruction_io_deq_bits_opcode == 4'h1 ? 3'h0 : _GEN_618; // @[Decoder.scala 282:51 669:15]
  assign lockPool_io_actor_1_out_ready = memPortBHandler_io_in_ready; // @[Decoder.scala 197:25]
  assign lockPool_io_lock_valid = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_46 : _GEN_601; // @[Decoder.scala 282:51]
  assign lockPool_io_lock_bits_cond_write = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_602; // @[Decoder.scala 282:51]
  assign lockPool_io_lock_bits_cond_address = instruction_io_deq_bits_opcode == 4'h1 ? args_memAddress : _GEN_603; // @[Decoder.scala 282:51]
  assign lockPool_io_lock_bits_cond_size = instruction_io_deq_bits_opcode == 4'h1 ? instruction_io_deq_ready_w_size :
    _GEN_604; // @[Decoder.scala 282:51]
  assign lockPool_io_lock_bits_cond_stride = instruction_io_deq_bits_opcode == 4'h1 ? args_memStride : _GEN_605; // @[Decoder.scala 282:51]
  assign lockPool_io_lock_bits_cond_reverse = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _T_3; // @[Decoder.scala 282:51]
  assign lockPool_io_lock_bits_lock = instruction_io_deq_bits_opcode == 4'h1 ? instruction_io_deq_ready_w_6_lock :
    _GEN_607; // @[Decoder.scala 282:51]
  assign lockPool_io_lock_bits_by = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_609; // @[Decoder.scala 282:51]
  assign accHandler_clock = clock;
  assign accHandler_reset = reset;
  assign accHandler_io_in_valid = acc_io_deq_valid; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_instruction_op = acc_io_deq_bits_instruction_op; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_instruction_sourceLeft = acc_io_deq_bits_instruction_sourceLeft; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_instruction_sourceRight = acc_io_deq_bits_instruction_sourceRight; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_instruction_dest = acc_io_deq_bits_instruction_dest; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_address = acc_io_deq_bits_address; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_altAddress = acc_io_deq_bits_altAddress; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_read = acc_io_deq_bits_read; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_write = acc_io_deq_bits_write; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_accumulate = acc_io_deq_bits_accumulate; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_size = acc_io_deq_bits_size; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_stride = acc_io_deq_bits_stride; // @[Mem.scala 23:7]
  assign accHandler_io_in_bits_reverse = acc_io_deq_bits_reverse; // @[Mem.scala 23:7]
  assign accHandler_io_out_ready = io_acc_ready; // @[Decoder.scala 219:27]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_io_enq_valid = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_20 : _GEN_632; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_instruction_op = instruction_io_deq_bits_opcode == 4'h1 ? 4'h0 : _GEN_633; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_instruction_sourceLeft = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_634; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_instruction_sourceRight = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_635; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_instruction_dest = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_636; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_address = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_25 : _GEN_637; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_altAddress = instruction_io_deq_bits_opcode == 4'h1 ? 12'h0 : _GEN_638; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_read = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_639; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_write = instruction_io_deq_bits_opcode == 4'h1 | _GEN_640; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_accumulate = instruction_io_deq_bits_opcode == 4'h1 ? flags_accumulate : _GEN_641; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_size = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_30 : _GEN_642; // @[Decoder.scala 282:51]
  assign acc_io_enq_bits_stride = instruction_io_deq_bits_opcode == 4'h1 ? args_accStride : _GEN_643; // @[Decoder.scala 282:51]
  assign acc_io_deq_ready = accHandler_io_in_ready; // @[Mem.scala 23:7]
  assign arrayHandler_clock = clock;
  assign arrayHandler_reset = reset;
  assign arrayHandler_io_in_valid = array_io_deq_valid; // @[Mem.scala 23:7]
  assign arrayHandler_io_in_bits_load = array_io_deq_bits_load; // @[Mem.scala 23:7]
  assign arrayHandler_io_in_bits_zeroes = array_io_deq_bits_zeroes; // @[Mem.scala 23:7]
  assign arrayHandler_io_in_bits_size = array_io_deq_bits_size; // @[Mem.scala 23:7]
  assign arrayHandler_io_out_ready = io_array_ready; // @[Decoder.scala 239:12]
  assign array_clock = clock;
  assign array_reset = reset;
  assign array_io_enq_valid = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_15 : _GEN_582; // @[Decoder.scala 282:51]
  assign array_io_enq_bits_load = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _T_3; // @[Decoder.scala 282:51]
  assign array_io_enq_bits_zeroes = instruction_io_deq_bits_opcode == 4'h1 ? flags_zeroes : _GEN_584; // @[Decoder.scala 282:51]
  assign array_io_enq_bits_size = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_13 : _GEN_585; // @[Decoder.scala 282:51]
  assign array_io_deq_ready = arrayHandler_io_in_ready; // @[Mem.scala 23:7]
  assign dataflow_clock = clock;
  assign dataflow_reset = reset;
  assign dataflow_io_enq_valid = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_11 : _GEN_589; // @[Decoder.scala 282:51]
  assign dataflow_io_enq_bits_kind = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_12 : _GEN_590; // @[Decoder.scala 282:51]
  assign dataflow_io_enq_bits_size = instruction_io_deq_bits_opcode == 4'h1 ? _GEN_13 : _GEN_591; // @[Decoder.scala 282:51]
  assign dataflow_io_deq_ready = io_dataflow_ready; // @[Mem.scala 23:7]
  assign hostDataflowHandler_clock = clock;
  assign hostDataflowHandler_reset = reset;
  assign hostDataflowHandler_io_in_valid = hostDataflow_io_deq_valid; // @[Mem.scala 23:7]
  assign hostDataflowHandler_io_in_bits_kind = hostDataflow_io_deq_bits_kind; // @[Mem.scala 23:7]
  assign hostDataflowHandler_io_in_bits_size = hostDataflow_io_deq_bits_size; // @[Mem.scala 23:7]
  assign hostDataflowHandler_io_out_ready = io_hostDataflow_ready; // @[Decoder.scala 257:19]
  assign hostDataflow_clock = clock;
  assign hostDataflow_reset = reset;
  assign hostDataflow_io_enq_valid = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_611; // @[Decoder.scala 282:51 670:16]
  assign hostDataflow_io_enq_bits_kind = instruction_io_deq_bits_opcode == 4'h1 ? 2'h0 : _GEN_612; // @[Decoder.scala 282:51 669:15]
  assign hostDataflow_io_enq_bits_size = instruction_io_deq_bits_opcode == 4'h1 ? 14'h0 : _GEN_613; // @[Decoder.scala 282:51 669:15]
  assign hostDataflow_io_deq_ready = hostDataflowHandler_io_in_ready; // @[Mem.scala 23:7]
  assign enqueuer1_clock = clock;
  assign enqueuer1_reset = reset;
  assign enqueuer1_io_in_valid = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_580; // @[Decoder.scala 282:51 MultiEnqueue.scala 40:17]
  assign enqueuer1_io_out_0_ready = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_581; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer2_clock = clock;
  assign enqueuer2_reset = reset;
  assign enqueuer2_io_in_valid = 1'h0; // @[MultiEnqueue.scala 40:17]
  assign enqueuer2_io_out_0_ready = 1'h0; // @[MultiEnqueue.scala 42:18]
  assign enqueuer2_io_out_1_ready = 1'h0; // @[MultiEnqueue.scala 42:18]
  assign enqueuer3_clock = clock;
  assign enqueuer3_reset = reset;
  assign enqueuer3_io_in_valid = instruction_io_deq_bits_opcode == 4'h1 & _GEN_9; // @[Decoder.scala 282:51 MultiEnqueue.scala 40:17]
  assign enqueuer3_io_out_0_ready = instruction_io_deq_bits_opcode == 4'h1 & _GEN_10; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer3_io_out_1_ready = instruction_io_deq_bits_opcode == 4'h1 & _GEN_14; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer3_io_out_2_ready = instruction_io_deq_bits_opcode == 4'h1 & _GEN_19; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer4_clock = clock;
  assign enqueuer4_reset = reset;
  assign enqueuer4_io_in_valid = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_587; // @[Decoder.scala 282:51 MultiEnqueue.scala 40:17]
  assign enqueuer4_io_out_0_ready = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_588; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer4_io_out_1_ready = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_592; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer4_io_out_2_ready = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_593; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer4_io_out_3_ready = instruction_io_deq_bits_opcode == 4'h1 ? 1'h0 : _GEN_600; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer5_clock = clock;
  assign enqueuer5_reset = reset;
  assign enqueuer5_io_in_valid = instruction_io_deq_bits_opcode == 4'h1 & _GEN_34; // @[Decoder.scala 282:51 MultiEnqueue.scala 40:17]
  assign enqueuer5_io_out_0_ready = instruction_io_deq_bits_opcode == 4'h1 & _GEN_35; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer5_io_out_1_ready = instruction_io_deq_bits_opcode == 4'h1 & _GEN_36; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer5_io_out_2_ready = instruction_io_deq_bits_opcode == 4'h1 & _GEN_43; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer5_io_out_3_ready = instruction_io_deq_bits_opcode == 4'h1 & _GEN_44; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  assign enqueuer5_io_out_4_ready = instruction_io_deq_bits_opcode == 4'h1 & _GEN_45; // @[Decoder.scala 282:51 MultiEnqueue.scala 42:18]
  always @(posedge clock) begin
    timeout <= _GEN_86[15:0]; // @[Decoder.scala 96:{24,24}]
    if (reset) begin // @[Decoder.scala 97:24]
      timer <= 16'h0; // @[Decoder.scala 97:24]
    end else if (instruction_io_deq_ready) begin // @[Decoder.scala 98:27]
      timer <= 16'h0; // @[Decoder.scala 99:11]
    end else if (timer < timeout) begin // @[Decoder.scala 101:27]
      timer <= _timer_T_1; // @[Decoder.scala 102:13]
    end
    if (reset) begin // @[Decoder.scala 108:31]
      tracepoint <= 32'hffffffff; // @[Decoder.scala 108:31]
    end else if (!(instruction_io_deq_bits_opcode == 4'h1)) begin // @[Decoder.scala 282:51]
      if (!(instruction_io_deq_bits_opcode == 4'h3)) begin // @[Decoder.scala 333:62]
        if (!(instruction_io_deq_bits_opcode == 4'h2)) begin // @[Decoder.scala 373:59]
          tracepoint <= _GEN_504;
        end
      end
    end
    if (reset) begin // @[Decoder.scala 109:31]
      programCounter <= 32'h0; // @[Decoder.scala 109:31]
    end else if (instruction_io_deq_bits_opcode == 4'h1) begin // @[Decoder.scala 282:51]
      programCounter <= _GEN_2;
    end else if (instruction_io_deq_bits_opcode == 4'h3) begin // @[Decoder.scala 333:62]
      programCounter <= _GEN_2;
    end else if (instruction_io_deq_bits_opcode == 4'h2) begin // @[Decoder.scala 373:59]
      programCounter <= _GEN_2;
    end else begin
      programCounter <= _GEN_505;
    end
    dram0AddressOffset <= _GEN_123[31:0]; // @[Decoder.scala 126:{35,35}]
    dram0CacheBehaviour <= _GEN_161[3:0]; // @[Decoder.scala 129:{36,36}]
    dram1AddressOffset <= _GEN_199[31:0]; // @[Decoder.scala 130:{35,35}]
    dram1CacheBehaviour <= _GEN_230[3:0]; // @[Decoder.scala 133:{36,36}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  timeout = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  timer = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  tracepoint = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  programCounter = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  dram0AddressOffset = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  dram0CacheBehaviour = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  dram1AddressOffset = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  dram1CacheBehaviour = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAC(
  input         clock,
  input         reset,
  input         io_load,
  input  [15:0] io_mulInput,
  input  [15:0] io_addInput,
  output [15:0] io_output,
  output [15:0] io_passthrough
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] weight; // @[MAC.scala 18:28]
  reg [15:0] passthrough; // @[MAC.scala 19:28]
  reg [24:0] output_; // @[MAC.scala 20:28]
  wire [31:0] _output_mac_T = $signed(io_mulInput) * $signed(weight); // @[package.scala 117:18]
  wire [23:0] _output_mac_T_1 = {$signed(io_addInput), 8'h0}; // @[package.scala 117:29]
  wire [31:0] _GEN_3 = {{8{_output_mac_T_1[23]}},_output_mac_T_1}; // @[package.scala 117:23]
  wire [32:0] output_mac = $signed(_output_mac_T) + $signed(_GEN_3); // @[package.scala 117:23]
  wire [8:0] output_mask1 = 9'sh80 - 9'sh1; // @[package.scala 120:44]
  wire [32:0] _output_adjustment_T_1 = $signed(output_mac) & 33'sh80; // @[package.scala 125:16]
  wire [32:0] _GEN_4 = {{24{output_mask1[8]}},output_mask1}; // @[package.scala 125:44]
  wire [32:0] _output_adjustment_T_4 = $signed(output_mac) & $signed(_GEN_4); // @[package.scala 125:44]
  wire [32:0] _output_adjustment_T_7 = $signed(output_mac) & 33'sh100; // @[package.scala 125:71]
  wire  _output_adjustment_T_10 = $signed(_output_adjustment_T_1) != 33'sh0 & ($signed(_output_adjustment_T_4) != 33'sh0
     | $signed(_output_adjustment_T_7) != 33'sh0); // @[package.scala 125:34]
  wire [1:0] output_adjustment = _output_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [24:0] _output_adjusted_T = output_mac[32:8]; // @[package.scala 130:26]
  wire [24:0] _GEN_5 = {{23{output_adjustment[1]}},output_adjustment}; // @[package.scala 130:42]
  wire [24:0] output_adjusted = $signed(_output_adjusted_T) + $signed(_GEN_5); // @[package.scala 130:42]
  wire [24:0] _GEN_1 = io_load ? $signed({{9{weight[15]}},weight}) : $signed(output_); // @[MAC.scala 25:17 27:15 30:15]
  assign io_output = _GEN_1[15:0];
  assign io_passthrough = passthrough; // @[MAC.scala 22:18]
  always @(posedge clock) begin
    if (reset) begin // @[MAC.scala 18:28]
      weight <= 16'sh0; // @[MAC.scala 18:28]
    end else if (io_load) begin // @[MAC.scala 25:17]
      weight <= io_addInput; // @[MAC.scala 26:12]
    end
    if (reset) begin // @[MAC.scala 19:28]
      passthrough <= 16'sh0; // @[MAC.scala 19:28]
    end else begin
      passthrough <= io_mulInput; // @[MAC.scala 23:15]
    end
    if (reset) begin // @[MAC.scala 20:28]
      output_ <= 25'sh0; // @[MAC.scala 20:28]
    end else if (!(io_load)) begin // @[MAC.scala 25:17]
      if ($signed(output_adjusted) > 25'sh7fff) begin // @[package.scala 98:8]
        output_ <= 25'sh7fff;
      end else if ($signed(output_adjusted) < -25'sh8000) begin // @[package.scala 98:26]
        output_ <= -25'sh8000;
      end else begin
        output_ <= output_adjusted;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  weight = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  passthrough = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  output_ = _RAND_2[24:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InnerSystolicArray(
  input         clock,
  input         reset,
  input         io_load,
  input  [15:0] io_input_0,
  input  [15:0] io_input_1,
  input  [15:0] io_input_2,
  input  [15:0] io_input_3,
  input  [15:0] io_input_4,
  input  [15:0] io_input_5,
  input  [15:0] io_input_6,
  input  [15:0] io_input_7,
  input  [15:0] io_input_8,
  input  [15:0] io_input_9,
  input  [15:0] io_input_10,
  input  [15:0] io_input_11,
  input  [15:0] io_input_12,
  input  [15:0] io_input_13,
  input  [15:0] io_input_14,
  input  [15:0] io_input_15,
  input  [15:0] io_input_16,
  input  [15:0] io_input_17,
  input  [15:0] io_input_18,
  input  [15:0] io_input_19,
  input  [15:0] io_input_20,
  input  [15:0] io_input_21,
  input  [15:0] io_input_22,
  input  [15:0] io_input_23,
  input  [15:0] io_input_24,
  input  [15:0] io_input_25,
  input  [15:0] io_input_26,
  input  [15:0] io_input_27,
  input  [15:0] io_input_28,
  input  [15:0] io_input_29,
  input  [15:0] io_input_30,
  input  [15:0] io_input_31,
  input  [15:0] io_weight_0,
  input  [15:0] io_weight_1,
  input  [15:0] io_weight_2,
  input  [15:0] io_weight_3,
  input  [15:0] io_weight_4,
  input  [15:0] io_weight_5,
  input  [15:0] io_weight_6,
  input  [15:0] io_weight_7,
  input  [15:0] io_weight_8,
  input  [15:0] io_weight_9,
  input  [15:0] io_weight_10,
  input  [15:0] io_weight_11,
  input  [15:0] io_weight_12,
  input  [15:0] io_weight_13,
  input  [15:0] io_weight_14,
  input  [15:0] io_weight_15,
  input  [15:0] io_weight_16,
  input  [15:0] io_weight_17,
  input  [15:0] io_weight_18,
  input  [15:0] io_weight_19,
  input  [15:0] io_weight_20,
  input  [15:0] io_weight_21,
  input  [15:0] io_weight_22,
  input  [15:0] io_weight_23,
  input  [15:0] io_weight_24,
  input  [15:0] io_weight_25,
  input  [15:0] io_weight_26,
  input  [15:0] io_weight_27,
  input  [15:0] io_weight_28,
  input  [15:0] io_weight_29,
  input  [15:0] io_weight_30,
  input  [15:0] io_weight_31,
  output [15:0] io_output_0,
  output [15:0] io_output_1,
  output [15:0] io_output_2,
  output [15:0] io_output_3,
  output [15:0] io_output_4,
  output [15:0] io_output_5,
  output [15:0] io_output_6,
  output [15:0] io_output_7,
  output [15:0] io_output_8,
  output [15:0] io_output_9,
  output [15:0] io_output_10,
  output [15:0] io_output_11,
  output [15:0] io_output_12,
  output [15:0] io_output_13,
  output [15:0] io_output_14,
  output [15:0] io_output_15,
  output [15:0] io_output_16,
  output [15:0] io_output_17,
  output [15:0] io_output_18,
  output [15:0] io_output_19,
  output [15:0] io_output_20,
  output [15:0] io_output_21,
  output [15:0] io_output_22,
  output [15:0] io_output_23,
  output [15:0] io_output_24,
  output [15:0] io_output_25,
  output [15:0] io_output_26,
  output [15:0] io_output_27,
  output [15:0] io_output_28,
  output [15:0] io_output_29,
  output [15:0] io_output_30,
  output [15:0] io_output_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
`endif // RANDOMIZE_REG_INIT
  wire  mac_0_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_0_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_0_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_1_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_1_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_2_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_2_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_3_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_3_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_4_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_4_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_5_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_5_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_6_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_6_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_7_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_7_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_8_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_8_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_9_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_9_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_10_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_10_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_11_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_11_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_12_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_12_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_13_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_13_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_14_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_14_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_15_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_15_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_16_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_16_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_17_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_17_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_18_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_18_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_19_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_19_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_20_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_20_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_21_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_21_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_22_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_22_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_23_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_23_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_24_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_24_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_25_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_25_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_26_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_26_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_27_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_27_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_28_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_28_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_29_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_29_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_30_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_30_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_0_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_0_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_0_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_0_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_0_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_0_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_0_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_1_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_1_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_1_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_1_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_1_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_1_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_1_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_2_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_2_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_2_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_2_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_2_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_2_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_2_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_3_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_3_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_3_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_3_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_3_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_3_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_3_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_4_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_4_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_4_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_4_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_4_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_4_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_4_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_5_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_5_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_5_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_5_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_5_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_5_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_5_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_6_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_6_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_6_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_6_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_6_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_6_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_6_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_7_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_7_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_7_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_7_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_7_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_7_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_7_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_8_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_8_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_8_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_8_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_8_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_8_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_8_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_9_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_9_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_9_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_9_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_9_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_9_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_9_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_10_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_10_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_10_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_10_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_10_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_10_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_10_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_11_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_11_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_11_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_11_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_11_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_11_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_11_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_12_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_12_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_12_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_12_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_12_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_12_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_12_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_13_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_13_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_13_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_13_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_13_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_13_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_13_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_14_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_14_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_14_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_14_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_14_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_14_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_14_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_15_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_15_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_15_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_15_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_15_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_15_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_15_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_16_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_16_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_16_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_16_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_16_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_16_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_16_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_17_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_17_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_17_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_17_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_17_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_17_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_17_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_18_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_18_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_18_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_18_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_18_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_18_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_18_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_19_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_19_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_19_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_19_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_19_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_19_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_19_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_20_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_20_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_20_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_20_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_20_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_20_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_20_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_21_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_21_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_21_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_21_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_21_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_21_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_21_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_22_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_22_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_22_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_22_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_22_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_22_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_22_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_23_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_23_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_23_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_23_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_23_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_23_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_23_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_24_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_24_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_24_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_24_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_24_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_24_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_24_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_25_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_25_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_25_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_25_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_25_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_25_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_25_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_26_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_26_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_26_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_26_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_26_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_26_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_26_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_27_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_27_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_27_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_27_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_27_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_27_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_27_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_28_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_28_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_28_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_28_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_28_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_28_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_28_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_29_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_29_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_29_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_29_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_29_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_29_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_29_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_30_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_30_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_30_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_30_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_30_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_30_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_30_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_31_clock; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_31_reset; // @[InnerSystolicArray.scala 34:50]
  wire  mac_31_31_io_load; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_31_io_mulInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_31_io_addInput; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_31_io_output; // @[InnerSystolicArray.scala 34:50]
  wire [15:0] mac_31_31_io_passthrough; // @[InnerSystolicArray.scala 34:50]
  reg [15:0] bias_0; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_1; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_2; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_3; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_4; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_5; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_6; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_7; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_8; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_9; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_10; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_11; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_12; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_13; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_14; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_15; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_16; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_17; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_18; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_19; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_20; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_21; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_22; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_23; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_24; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_25; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_26; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_27; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_28; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_29; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_30; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] bias_31; // @[InnerSystolicArray.scala 37:20]
  reg [15:0] mac_0_1_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_2_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_2_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_3_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_3_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_3_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_4_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_4_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_4_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_4_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_5_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_5_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_5_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_5_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_5_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_6_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_6_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_6_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_6_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_6_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_6_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_7_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_7_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_7_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_7_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_7_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_7_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_7_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_8_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_8_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_8_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_8_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_8_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_8_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_8_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_8_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_9_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_9_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_9_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_9_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_9_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_9_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_9_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_9_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_9_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_10_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_10_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_10_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_10_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_10_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_10_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_10_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_10_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_10_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_10_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_11_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_12_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_13_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_14_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_15_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_16_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_17_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_18_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_19_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_20_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_21_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_22_io_mulInput_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_23_io_mulInput_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_24_io_mulInput_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_25_io_mulInput_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_26_io_mulInput_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_27_io_mulInput_sr_26; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_26; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_28_io_mulInput_sr_27; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_26; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_27; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_29_io_mulInput_sr_28; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_26; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_27; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_28; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_30_io_mulInput_sr_29; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_26; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_27; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_28; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_29; // @[ShiftRegister.scala 10:22]
  reg [15:0] mac_0_31_io_mulInput_sr_30; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_26; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_27; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_28; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_29; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_0_sr_30; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_26; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_27; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_28; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_1_sr_29; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_26; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_27; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_2_sr_28; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_26; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_3_sr_27; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_4_sr_26; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_5_sr_25; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_6_sr_24; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_7_sr_23; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_8_sr_22; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_9_sr_21; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_10_sr_20; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_11_sr_19; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_12_sr_18; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_13_sr_17; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_14_sr_16; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_15_sr_15; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_16_sr_14; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_17_sr_13; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_18_sr_12; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_19_sr_11; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_20_sr_10; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_21_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_21_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_21_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_21_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_21_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_21_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_21_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_21_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_21_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_21_sr_9; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_22_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_22_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_22_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_22_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_22_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_22_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_22_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_22_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_22_sr_8; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_23_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_23_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_23_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_23_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_23_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_23_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_23_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_23_sr_7; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_24_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_24_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_24_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_24_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_24_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_24_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_24_sr_6; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_25_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_25_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_25_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_25_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_25_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_25_sr_5; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_26_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_26_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_26_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_26_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_26_sr_4; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_27_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_27_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_27_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_27_sr_3; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_28_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_28_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_28_sr_2; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_29_sr_0; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_29_sr_1; // @[ShiftRegister.scala 10:22]
  reg [15:0] io_output_30_sr_0; // @[ShiftRegister.scala 10:22]
  MAC mac_0_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_0_clock),
    .reset(mac_0_0_reset),
    .io_load(mac_0_0_io_load),
    .io_mulInput(mac_0_0_io_mulInput),
    .io_addInput(mac_0_0_io_addInput),
    .io_output(mac_0_0_io_output),
    .io_passthrough(mac_0_0_io_passthrough)
  );
  MAC mac_0_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_1_clock),
    .reset(mac_0_1_reset),
    .io_load(mac_0_1_io_load),
    .io_mulInput(mac_0_1_io_mulInput),
    .io_addInput(mac_0_1_io_addInput),
    .io_output(mac_0_1_io_output),
    .io_passthrough(mac_0_1_io_passthrough)
  );
  MAC mac_0_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_2_clock),
    .reset(mac_0_2_reset),
    .io_load(mac_0_2_io_load),
    .io_mulInput(mac_0_2_io_mulInput),
    .io_addInput(mac_0_2_io_addInput),
    .io_output(mac_0_2_io_output),
    .io_passthrough(mac_0_2_io_passthrough)
  );
  MAC mac_0_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_3_clock),
    .reset(mac_0_3_reset),
    .io_load(mac_0_3_io_load),
    .io_mulInput(mac_0_3_io_mulInput),
    .io_addInput(mac_0_3_io_addInput),
    .io_output(mac_0_3_io_output),
    .io_passthrough(mac_0_3_io_passthrough)
  );
  MAC mac_0_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_4_clock),
    .reset(mac_0_4_reset),
    .io_load(mac_0_4_io_load),
    .io_mulInput(mac_0_4_io_mulInput),
    .io_addInput(mac_0_4_io_addInput),
    .io_output(mac_0_4_io_output),
    .io_passthrough(mac_0_4_io_passthrough)
  );
  MAC mac_0_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_5_clock),
    .reset(mac_0_5_reset),
    .io_load(mac_0_5_io_load),
    .io_mulInput(mac_0_5_io_mulInput),
    .io_addInput(mac_0_5_io_addInput),
    .io_output(mac_0_5_io_output),
    .io_passthrough(mac_0_5_io_passthrough)
  );
  MAC mac_0_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_6_clock),
    .reset(mac_0_6_reset),
    .io_load(mac_0_6_io_load),
    .io_mulInput(mac_0_6_io_mulInput),
    .io_addInput(mac_0_6_io_addInput),
    .io_output(mac_0_6_io_output),
    .io_passthrough(mac_0_6_io_passthrough)
  );
  MAC mac_0_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_7_clock),
    .reset(mac_0_7_reset),
    .io_load(mac_0_7_io_load),
    .io_mulInput(mac_0_7_io_mulInput),
    .io_addInput(mac_0_7_io_addInput),
    .io_output(mac_0_7_io_output),
    .io_passthrough(mac_0_7_io_passthrough)
  );
  MAC mac_0_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_8_clock),
    .reset(mac_0_8_reset),
    .io_load(mac_0_8_io_load),
    .io_mulInput(mac_0_8_io_mulInput),
    .io_addInput(mac_0_8_io_addInput),
    .io_output(mac_0_8_io_output),
    .io_passthrough(mac_0_8_io_passthrough)
  );
  MAC mac_0_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_9_clock),
    .reset(mac_0_9_reset),
    .io_load(mac_0_9_io_load),
    .io_mulInput(mac_0_9_io_mulInput),
    .io_addInput(mac_0_9_io_addInput),
    .io_output(mac_0_9_io_output),
    .io_passthrough(mac_0_9_io_passthrough)
  );
  MAC mac_0_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_10_clock),
    .reset(mac_0_10_reset),
    .io_load(mac_0_10_io_load),
    .io_mulInput(mac_0_10_io_mulInput),
    .io_addInput(mac_0_10_io_addInput),
    .io_output(mac_0_10_io_output),
    .io_passthrough(mac_0_10_io_passthrough)
  );
  MAC mac_0_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_11_clock),
    .reset(mac_0_11_reset),
    .io_load(mac_0_11_io_load),
    .io_mulInput(mac_0_11_io_mulInput),
    .io_addInput(mac_0_11_io_addInput),
    .io_output(mac_0_11_io_output),
    .io_passthrough(mac_0_11_io_passthrough)
  );
  MAC mac_0_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_12_clock),
    .reset(mac_0_12_reset),
    .io_load(mac_0_12_io_load),
    .io_mulInput(mac_0_12_io_mulInput),
    .io_addInput(mac_0_12_io_addInput),
    .io_output(mac_0_12_io_output),
    .io_passthrough(mac_0_12_io_passthrough)
  );
  MAC mac_0_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_13_clock),
    .reset(mac_0_13_reset),
    .io_load(mac_0_13_io_load),
    .io_mulInput(mac_0_13_io_mulInput),
    .io_addInput(mac_0_13_io_addInput),
    .io_output(mac_0_13_io_output),
    .io_passthrough(mac_0_13_io_passthrough)
  );
  MAC mac_0_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_14_clock),
    .reset(mac_0_14_reset),
    .io_load(mac_0_14_io_load),
    .io_mulInput(mac_0_14_io_mulInput),
    .io_addInput(mac_0_14_io_addInput),
    .io_output(mac_0_14_io_output),
    .io_passthrough(mac_0_14_io_passthrough)
  );
  MAC mac_0_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_15_clock),
    .reset(mac_0_15_reset),
    .io_load(mac_0_15_io_load),
    .io_mulInput(mac_0_15_io_mulInput),
    .io_addInput(mac_0_15_io_addInput),
    .io_output(mac_0_15_io_output),
    .io_passthrough(mac_0_15_io_passthrough)
  );
  MAC mac_0_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_16_clock),
    .reset(mac_0_16_reset),
    .io_load(mac_0_16_io_load),
    .io_mulInput(mac_0_16_io_mulInput),
    .io_addInput(mac_0_16_io_addInput),
    .io_output(mac_0_16_io_output),
    .io_passthrough(mac_0_16_io_passthrough)
  );
  MAC mac_0_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_17_clock),
    .reset(mac_0_17_reset),
    .io_load(mac_0_17_io_load),
    .io_mulInput(mac_0_17_io_mulInput),
    .io_addInput(mac_0_17_io_addInput),
    .io_output(mac_0_17_io_output),
    .io_passthrough(mac_0_17_io_passthrough)
  );
  MAC mac_0_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_18_clock),
    .reset(mac_0_18_reset),
    .io_load(mac_0_18_io_load),
    .io_mulInput(mac_0_18_io_mulInput),
    .io_addInput(mac_0_18_io_addInput),
    .io_output(mac_0_18_io_output),
    .io_passthrough(mac_0_18_io_passthrough)
  );
  MAC mac_0_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_19_clock),
    .reset(mac_0_19_reset),
    .io_load(mac_0_19_io_load),
    .io_mulInput(mac_0_19_io_mulInput),
    .io_addInput(mac_0_19_io_addInput),
    .io_output(mac_0_19_io_output),
    .io_passthrough(mac_0_19_io_passthrough)
  );
  MAC mac_0_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_20_clock),
    .reset(mac_0_20_reset),
    .io_load(mac_0_20_io_load),
    .io_mulInput(mac_0_20_io_mulInput),
    .io_addInput(mac_0_20_io_addInput),
    .io_output(mac_0_20_io_output),
    .io_passthrough(mac_0_20_io_passthrough)
  );
  MAC mac_0_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_21_clock),
    .reset(mac_0_21_reset),
    .io_load(mac_0_21_io_load),
    .io_mulInput(mac_0_21_io_mulInput),
    .io_addInput(mac_0_21_io_addInput),
    .io_output(mac_0_21_io_output),
    .io_passthrough(mac_0_21_io_passthrough)
  );
  MAC mac_0_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_22_clock),
    .reset(mac_0_22_reset),
    .io_load(mac_0_22_io_load),
    .io_mulInput(mac_0_22_io_mulInput),
    .io_addInput(mac_0_22_io_addInput),
    .io_output(mac_0_22_io_output),
    .io_passthrough(mac_0_22_io_passthrough)
  );
  MAC mac_0_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_23_clock),
    .reset(mac_0_23_reset),
    .io_load(mac_0_23_io_load),
    .io_mulInput(mac_0_23_io_mulInput),
    .io_addInput(mac_0_23_io_addInput),
    .io_output(mac_0_23_io_output),
    .io_passthrough(mac_0_23_io_passthrough)
  );
  MAC mac_0_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_24_clock),
    .reset(mac_0_24_reset),
    .io_load(mac_0_24_io_load),
    .io_mulInput(mac_0_24_io_mulInput),
    .io_addInput(mac_0_24_io_addInput),
    .io_output(mac_0_24_io_output),
    .io_passthrough(mac_0_24_io_passthrough)
  );
  MAC mac_0_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_25_clock),
    .reset(mac_0_25_reset),
    .io_load(mac_0_25_io_load),
    .io_mulInput(mac_0_25_io_mulInput),
    .io_addInput(mac_0_25_io_addInput),
    .io_output(mac_0_25_io_output),
    .io_passthrough(mac_0_25_io_passthrough)
  );
  MAC mac_0_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_26_clock),
    .reset(mac_0_26_reset),
    .io_load(mac_0_26_io_load),
    .io_mulInput(mac_0_26_io_mulInput),
    .io_addInput(mac_0_26_io_addInput),
    .io_output(mac_0_26_io_output),
    .io_passthrough(mac_0_26_io_passthrough)
  );
  MAC mac_0_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_27_clock),
    .reset(mac_0_27_reset),
    .io_load(mac_0_27_io_load),
    .io_mulInput(mac_0_27_io_mulInput),
    .io_addInput(mac_0_27_io_addInput),
    .io_output(mac_0_27_io_output),
    .io_passthrough(mac_0_27_io_passthrough)
  );
  MAC mac_0_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_28_clock),
    .reset(mac_0_28_reset),
    .io_load(mac_0_28_io_load),
    .io_mulInput(mac_0_28_io_mulInput),
    .io_addInput(mac_0_28_io_addInput),
    .io_output(mac_0_28_io_output),
    .io_passthrough(mac_0_28_io_passthrough)
  );
  MAC mac_0_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_29_clock),
    .reset(mac_0_29_reset),
    .io_load(mac_0_29_io_load),
    .io_mulInput(mac_0_29_io_mulInput),
    .io_addInput(mac_0_29_io_addInput),
    .io_output(mac_0_29_io_output),
    .io_passthrough(mac_0_29_io_passthrough)
  );
  MAC mac_0_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_30_clock),
    .reset(mac_0_30_reset),
    .io_load(mac_0_30_io_load),
    .io_mulInput(mac_0_30_io_mulInput),
    .io_addInput(mac_0_30_io_addInput),
    .io_output(mac_0_30_io_output),
    .io_passthrough(mac_0_30_io_passthrough)
  );
  MAC mac_0_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_0_31_clock),
    .reset(mac_0_31_reset),
    .io_load(mac_0_31_io_load),
    .io_mulInput(mac_0_31_io_mulInput),
    .io_addInput(mac_0_31_io_addInput),
    .io_output(mac_0_31_io_output),
    .io_passthrough(mac_0_31_io_passthrough)
  );
  MAC mac_1_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_0_clock),
    .reset(mac_1_0_reset),
    .io_load(mac_1_0_io_load),
    .io_mulInput(mac_1_0_io_mulInput),
    .io_addInput(mac_1_0_io_addInput),
    .io_output(mac_1_0_io_output),
    .io_passthrough(mac_1_0_io_passthrough)
  );
  MAC mac_1_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_1_clock),
    .reset(mac_1_1_reset),
    .io_load(mac_1_1_io_load),
    .io_mulInput(mac_1_1_io_mulInput),
    .io_addInput(mac_1_1_io_addInput),
    .io_output(mac_1_1_io_output),
    .io_passthrough(mac_1_1_io_passthrough)
  );
  MAC mac_1_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_2_clock),
    .reset(mac_1_2_reset),
    .io_load(mac_1_2_io_load),
    .io_mulInput(mac_1_2_io_mulInput),
    .io_addInput(mac_1_2_io_addInput),
    .io_output(mac_1_2_io_output),
    .io_passthrough(mac_1_2_io_passthrough)
  );
  MAC mac_1_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_3_clock),
    .reset(mac_1_3_reset),
    .io_load(mac_1_3_io_load),
    .io_mulInput(mac_1_3_io_mulInput),
    .io_addInput(mac_1_3_io_addInput),
    .io_output(mac_1_3_io_output),
    .io_passthrough(mac_1_3_io_passthrough)
  );
  MAC mac_1_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_4_clock),
    .reset(mac_1_4_reset),
    .io_load(mac_1_4_io_load),
    .io_mulInput(mac_1_4_io_mulInput),
    .io_addInput(mac_1_4_io_addInput),
    .io_output(mac_1_4_io_output),
    .io_passthrough(mac_1_4_io_passthrough)
  );
  MAC mac_1_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_5_clock),
    .reset(mac_1_5_reset),
    .io_load(mac_1_5_io_load),
    .io_mulInput(mac_1_5_io_mulInput),
    .io_addInput(mac_1_5_io_addInput),
    .io_output(mac_1_5_io_output),
    .io_passthrough(mac_1_5_io_passthrough)
  );
  MAC mac_1_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_6_clock),
    .reset(mac_1_6_reset),
    .io_load(mac_1_6_io_load),
    .io_mulInput(mac_1_6_io_mulInput),
    .io_addInput(mac_1_6_io_addInput),
    .io_output(mac_1_6_io_output),
    .io_passthrough(mac_1_6_io_passthrough)
  );
  MAC mac_1_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_7_clock),
    .reset(mac_1_7_reset),
    .io_load(mac_1_7_io_load),
    .io_mulInput(mac_1_7_io_mulInput),
    .io_addInput(mac_1_7_io_addInput),
    .io_output(mac_1_7_io_output),
    .io_passthrough(mac_1_7_io_passthrough)
  );
  MAC mac_1_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_8_clock),
    .reset(mac_1_8_reset),
    .io_load(mac_1_8_io_load),
    .io_mulInput(mac_1_8_io_mulInput),
    .io_addInput(mac_1_8_io_addInput),
    .io_output(mac_1_8_io_output),
    .io_passthrough(mac_1_8_io_passthrough)
  );
  MAC mac_1_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_9_clock),
    .reset(mac_1_9_reset),
    .io_load(mac_1_9_io_load),
    .io_mulInput(mac_1_9_io_mulInput),
    .io_addInput(mac_1_9_io_addInput),
    .io_output(mac_1_9_io_output),
    .io_passthrough(mac_1_9_io_passthrough)
  );
  MAC mac_1_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_10_clock),
    .reset(mac_1_10_reset),
    .io_load(mac_1_10_io_load),
    .io_mulInput(mac_1_10_io_mulInput),
    .io_addInput(mac_1_10_io_addInput),
    .io_output(mac_1_10_io_output),
    .io_passthrough(mac_1_10_io_passthrough)
  );
  MAC mac_1_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_11_clock),
    .reset(mac_1_11_reset),
    .io_load(mac_1_11_io_load),
    .io_mulInput(mac_1_11_io_mulInput),
    .io_addInput(mac_1_11_io_addInput),
    .io_output(mac_1_11_io_output),
    .io_passthrough(mac_1_11_io_passthrough)
  );
  MAC mac_1_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_12_clock),
    .reset(mac_1_12_reset),
    .io_load(mac_1_12_io_load),
    .io_mulInput(mac_1_12_io_mulInput),
    .io_addInput(mac_1_12_io_addInput),
    .io_output(mac_1_12_io_output),
    .io_passthrough(mac_1_12_io_passthrough)
  );
  MAC mac_1_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_13_clock),
    .reset(mac_1_13_reset),
    .io_load(mac_1_13_io_load),
    .io_mulInput(mac_1_13_io_mulInput),
    .io_addInput(mac_1_13_io_addInput),
    .io_output(mac_1_13_io_output),
    .io_passthrough(mac_1_13_io_passthrough)
  );
  MAC mac_1_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_14_clock),
    .reset(mac_1_14_reset),
    .io_load(mac_1_14_io_load),
    .io_mulInput(mac_1_14_io_mulInput),
    .io_addInput(mac_1_14_io_addInput),
    .io_output(mac_1_14_io_output),
    .io_passthrough(mac_1_14_io_passthrough)
  );
  MAC mac_1_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_15_clock),
    .reset(mac_1_15_reset),
    .io_load(mac_1_15_io_load),
    .io_mulInput(mac_1_15_io_mulInput),
    .io_addInput(mac_1_15_io_addInput),
    .io_output(mac_1_15_io_output),
    .io_passthrough(mac_1_15_io_passthrough)
  );
  MAC mac_1_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_16_clock),
    .reset(mac_1_16_reset),
    .io_load(mac_1_16_io_load),
    .io_mulInput(mac_1_16_io_mulInput),
    .io_addInput(mac_1_16_io_addInput),
    .io_output(mac_1_16_io_output),
    .io_passthrough(mac_1_16_io_passthrough)
  );
  MAC mac_1_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_17_clock),
    .reset(mac_1_17_reset),
    .io_load(mac_1_17_io_load),
    .io_mulInput(mac_1_17_io_mulInput),
    .io_addInput(mac_1_17_io_addInput),
    .io_output(mac_1_17_io_output),
    .io_passthrough(mac_1_17_io_passthrough)
  );
  MAC mac_1_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_18_clock),
    .reset(mac_1_18_reset),
    .io_load(mac_1_18_io_load),
    .io_mulInput(mac_1_18_io_mulInput),
    .io_addInput(mac_1_18_io_addInput),
    .io_output(mac_1_18_io_output),
    .io_passthrough(mac_1_18_io_passthrough)
  );
  MAC mac_1_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_19_clock),
    .reset(mac_1_19_reset),
    .io_load(mac_1_19_io_load),
    .io_mulInput(mac_1_19_io_mulInput),
    .io_addInput(mac_1_19_io_addInput),
    .io_output(mac_1_19_io_output),
    .io_passthrough(mac_1_19_io_passthrough)
  );
  MAC mac_1_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_20_clock),
    .reset(mac_1_20_reset),
    .io_load(mac_1_20_io_load),
    .io_mulInput(mac_1_20_io_mulInput),
    .io_addInput(mac_1_20_io_addInput),
    .io_output(mac_1_20_io_output),
    .io_passthrough(mac_1_20_io_passthrough)
  );
  MAC mac_1_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_21_clock),
    .reset(mac_1_21_reset),
    .io_load(mac_1_21_io_load),
    .io_mulInput(mac_1_21_io_mulInput),
    .io_addInput(mac_1_21_io_addInput),
    .io_output(mac_1_21_io_output),
    .io_passthrough(mac_1_21_io_passthrough)
  );
  MAC mac_1_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_22_clock),
    .reset(mac_1_22_reset),
    .io_load(mac_1_22_io_load),
    .io_mulInput(mac_1_22_io_mulInput),
    .io_addInput(mac_1_22_io_addInput),
    .io_output(mac_1_22_io_output),
    .io_passthrough(mac_1_22_io_passthrough)
  );
  MAC mac_1_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_23_clock),
    .reset(mac_1_23_reset),
    .io_load(mac_1_23_io_load),
    .io_mulInput(mac_1_23_io_mulInput),
    .io_addInput(mac_1_23_io_addInput),
    .io_output(mac_1_23_io_output),
    .io_passthrough(mac_1_23_io_passthrough)
  );
  MAC mac_1_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_24_clock),
    .reset(mac_1_24_reset),
    .io_load(mac_1_24_io_load),
    .io_mulInput(mac_1_24_io_mulInput),
    .io_addInput(mac_1_24_io_addInput),
    .io_output(mac_1_24_io_output),
    .io_passthrough(mac_1_24_io_passthrough)
  );
  MAC mac_1_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_25_clock),
    .reset(mac_1_25_reset),
    .io_load(mac_1_25_io_load),
    .io_mulInput(mac_1_25_io_mulInput),
    .io_addInput(mac_1_25_io_addInput),
    .io_output(mac_1_25_io_output),
    .io_passthrough(mac_1_25_io_passthrough)
  );
  MAC mac_1_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_26_clock),
    .reset(mac_1_26_reset),
    .io_load(mac_1_26_io_load),
    .io_mulInput(mac_1_26_io_mulInput),
    .io_addInput(mac_1_26_io_addInput),
    .io_output(mac_1_26_io_output),
    .io_passthrough(mac_1_26_io_passthrough)
  );
  MAC mac_1_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_27_clock),
    .reset(mac_1_27_reset),
    .io_load(mac_1_27_io_load),
    .io_mulInput(mac_1_27_io_mulInput),
    .io_addInput(mac_1_27_io_addInput),
    .io_output(mac_1_27_io_output),
    .io_passthrough(mac_1_27_io_passthrough)
  );
  MAC mac_1_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_28_clock),
    .reset(mac_1_28_reset),
    .io_load(mac_1_28_io_load),
    .io_mulInput(mac_1_28_io_mulInput),
    .io_addInput(mac_1_28_io_addInput),
    .io_output(mac_1_28_io_output),
    .io_passthrough(mac_1_28_io_passthrough)
  );
  MAC mac_1_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_29_clock),
    .reset(mac_1_29_reset),
    .io_load(mac_1_29_io_load),
    .io_mulInput(mac_1_29_io_mulInput),
    .io_addInput(mac_1_29_io_addInput),
    .io_output(mac_1_29_io_output),
    .io_passthrough(mac_1_29_io_passthrough)
  );
  MAC mac_1_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_30_clock),
    .reset(mac_1_30_reset),
    .io_load(mac_1_30_io_load),
    .io_mulInput(mac_1_30_io_mulInput),
    .io_addInput(mac_1_30_io_addInput),
    .io_output(mac_1_30_io_output),
    .io_passthrough(mac_1_30_io_passthrough)
  );
  MAC mac_1_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_1_31_clock),
    .reset(mac_1_31_reset),
    .io_load(mac_1_31_io_load),
    .io_mulInput(mac_1_31_io_mulInput),
    .io_addInput(mac_1_31_io_addInput),
    .io_output(mac_1_31_io_output),
    .io_passthrough(mac_1_31_io_passthrough)
  );
  MAC mac_2_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_0_clock),
    .reset(mac_2_0_reset),
    .io_load(mac_2_0_io_load),
    .io_mulInput(mac_2_0_io_mulInput),
    .io_addInput(mac_2_0_io_addInput),
    .io_output(mac_2_0_io_output),
    .io_passthrough(mac_2_0_io_passthrough)
  );
  MAC mac_2_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_1_clock),
    .reset(mac_2_1_reset),
    .io_load(mac_2_1_io_load),
    .io_mulInput(mac_2_1_io_mulInput),
    .io_addInput(mac_2_1_io_addInput),
    .io_output(mac_2_1_io_output),
    .io_passthrough(mac_2_1_io_passthrough)
  );
  MAC mac_2_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_2_clock),
    .reset(mac_2_2_reset),
    .io_load(mac_2_2_io_load),
    .io_mulInput(mac_2_2_io_mulInput),
    .io_addInput(mac_2_2_io_addInput),
    .io_output(mac_2_2_io_output),
    .io_passthrough(mac_2_2_io_passthrough)
  );
  MAC mac_2_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_3_clock),
    .reset(mac_2_3_reset),
    .io_load(mac_2_3_io_load),
    .io_mulInput(mac_2_3_io_mulInput),
    .io_addInput(mac_2_3_io_addInput),
    .io_output(mac_2_3_io_output),
    .io_passthrough(mac_2_3_io_passthrough)
  );
  MAC mac_2_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_4_clock),
    .reset(mac_2_4_reset),
    .io_load(mac_2_4_io_load),
    .io_mulInput(mac_2_4_io_mulInput),
    .io_addInput(mac_2_4_io_addInput),
    .io_output(mac_2_4_io_output),
    .io_passthrough(mac_2_4_io_passthrough)
  );
  MAC mac_2_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_5_clock),
    .reset(mac_2_5_reset),
    .io_load(mac_2_5_io_load),
    .io_mulInput(mac_2_5_io_mulInput),
    .io_addInput(mac_2_5_io_addInput),
    .io_output(mac_2_5_io_output),
    .io_passthrough(mac_2_5_io_passthrough)
  );
  MAC mac_2_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_6_clock),
    .reset(mac_2_6_reset),
    .io_load(mac_2_6_io_load),
    .io_mulInput(mac_2_6_io_mulInput),
    .io_addInput(mac_2_6_io_addInput),
    .io_output(mac_2_6_io_output),
    .io_passthrough(mac_2_6_io_passthrough)
  );
  MAC mac_2_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_7_clock),
    .reset(mac_2_7_reset),
    .io_load(mac_2_7_io_load),
    .io_mulInput(mac_2_7_io_mulInput),
    .io_addInput(mac_2_7_io_addInput),
    .io_output(mac_2_7_io_output),
    .io_passthrough(mac_2_7_io_passthrough)
  );
  MAC mac_2_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_8_clock),
    .reset(mac_2_8_reset),
    .io_load(mac_2_8_io_load),
    .io_mulInput(mac_2_8_io_mulInput),
    .io_addInput(mac_2_8_io_addInput),
    .io_output(mac_2_8_io_output),
    .io_passthrough(mac_2_8_io_passthrough)
  );
  MAC mac_2_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_9_clock),
    .reset(mac_2_9_reset),
    .io_load(mac_2_9_io_load),
    .io_mulInput(mac_2_9_io_mulInput),
    .io_addInput(mac_2_9_io_addInput),
    .io_output(mac_2_9_io_output),
    .io_passthrough(mac_2_9_io_passthrough)
  );
  MAC mac_2_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_10_clock),
    .reset(mac_2_10_reset),
    .io_load(mac_2_10_io_load),
    .io_mulInput(mac_2_10_io_mulInput),
    .io_addInput(mac_2_10_io_addInput),
    .io_output(mac_2_10_io_output),
    .io_passthrough(mac_2_10_io_passthrough)
  );
  MAC mac_2_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_11_clock),
    .reset(mac_2_11_reset),
    .io_load(mac_2_11_io_load),
    .io_mulInput(mac_2_11_io_mulInput),
    .io_addInput(mac_2_11_io_addInput),
    .io_output(mac_2_11_io_output),
    .io_passthrough(mac_2_11_io_passthrough)
  );
  MAC mac_2_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_12_clock),
    .reset(mac_2_12_reset),
    .io_load(mac_2_12_io_load),
    .io_mulInput(mac_2_12_io_mulInput),
    .io_addInput(mac_2_12_io_addInput),
    .io_output(mac_2_12_io_output),
    .io_passthrough(mac_2_12_io_passthrough)
  );
  MAC mac_2_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_13_clock),
    .reset(mac_2_13_reset),
    .io_load(mac_2_13_io_load),
    .io_mulInput(mac_2_13_io_mulInput),
    .io_addInput(mac_2_13_io_addInput),
    .io_output(mac_2_13_io_output),
    .io_passthrough(mac_2_13_io_passthrough)
  );
  MAC mac_2_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_14_clock),
    .reset(mac_2_14_reset),
    .io_load(mac_2_14_io_load),
    .io_mulInput(mac_2_14_io_mulInput),
    .io_addInput(mac_2_14_io_addInput),
    .io_output(mac_2_14_io_output),
    .io_passthrough(mac_2_14_io_passthrough)
  );
  MAC mac_2_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_15_clock),
    .reset(mac_2_15_reset),
    .io_load(mac_2_15_io_load),
    .io_mulInput(mac_2_15_io_mulInput),
    .io_addInput(mac_2_15_io_addInput),
    .io_output(mac_2_15_io_output),
    .io_passthrough(mac_2_15_io_passthrough)
  );
  MAC mac_2_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_16_clock),
    .reset(mac_2_16_reset),
    .io_load(mac_2_16_io_load),
    .io_mulInput(mac_2_16_io_mulInput),
    .io_addInput(mac_2_16_io_addInput),
    .io_output(mac_2_16_io_output),
    .io_passthrough(mac_2_16_io_passthrough)
  );
  MAC mac_2_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_17_clock),
    .reset(mac_2_17_reset),
    .io_load(mac_2_17_io_load),
    .io_mulInput(mac_2_17_io_mulInput),
    .io_addInput(mac_2_17_io_addInput),
    .io_output(mac_2_17_io_output),
    .io_passthrough(mac_2_17_io_passthrough)
  );
  MAC mac_2_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_18_clock),
    .reset(mac_2_18_reset),
    .io_load(mac_2_18_io_load),
    .io_mulInput(mac_2_18_io_mulInput),
    .io_addInput(mac_2_18_io_addInput),
    .io_output(mac_2_18_io_output),
    .io_passthrough(mac_2_18_io_passthrough)
  );
  MAC mac_2_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_19_clock),
    .reset(mac_2_19_reset),
    .io_load(mac_2_19_io_load),
    .io_mulInput(mac_2_19_io_mulInput),
    .io_addInput(mac_2_19_io_addInput),
    .io_output(mac_2_19_io_output),
    .io_passthrough(mac_2_19_io_passthrough)
  );
  MAC mac_2_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_20_clock),
    .reset(mac_2_20_reset),
    .io_load(mac_2_20_io_load),
    .io_mulInput(mac_2_20_io_mulInput),
    .io_addInput(mac_2_20_io_addInput),
    .io_output(mac_2_20_io_output),
    .io_passthrough(mac_2_20_io_passthrough)
  );
  MAC mac_2_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_21_clock),
    .reset(mac_2_21_reset),
    .io_load(mac_2_21_io_load),
    .io_mulInput(mac_2_21_io_mulInput),
    .io_addInput(mac_2_21_io_addInput),
    .io_output(mac_2_21_io_output),
    .io_passthrough(mac_2_21_io_passthrough)
  );
  MAC mac_2_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_22_clock),
    .reset(mac_2_22_reset),
    .io_load(mac_2_22_io_load),
    .io_mulInput(mac_2_22_io_mulInput),
    .io_addInput(mac_2_22_io_addInput),
    .io_output(mac_2_22_io_output),
    .io_passthrough(mac_2_22_io_passthrough)
  );
  MAC mac_2_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_23_clock),
    .reset(mac_2_23_reset),
    .io_load(mac_2_23_io_load),
    .io_mulInput(mac_2_23_io_mulInput),
    .io_addInput(mac_2_23_io_addInput),
    .io_output(mac_2_23_io_output),
    .io_passthrough(mac_2_23_io_passthrough)
  );
  MAC mac_2_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_24_clock),
    .reset(mac_2_24_reset),
    .io_load(mac_2_24_io_load),
    .io_mulInput(mac_2_24_io_mulInput),
    .io_addInput(mac_2_24_io_addInput),
    .io_output(mac_2_24_io_output),
    .io_passthrough(mac_2_24_io_passthrough)
  );
  MAC mac_2_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_25_clock),
    .reset(mac_2_25_reset),
    .io_load(mac_2_25_io_load),
    .io_mulInput(mac_2_25_io_mulInput),
    .io_addInput(mac_2_25_io_addInput),
    .io_output(mac_2_25_io_output),
    .io_passthrough(mac_2_25_io_passthrough)
  );
  MAC mac_2_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_26_clock),
    .reset(mac_2_26_reset),
    .io_load(mac_2_26_io_load),
    .io_mulInput(mac_2_26_io_mulInput),
    .io_addInput(mac_2_26_io_addInput),
    .io_output(mac_2_26_io_output),
    .io_passthrough(mac_2_26_io_passthrough)
  );
  MAC mac_2_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_27_clock),
    .reset(mac_2_27_reset),
    .io_load(mac_2_27_io_load),
    .io_mulInput(mac_2_27_io_mulInput),
    .io_addInput(mac_2_27_io_addInput),
    .io_output(mac_2_27_io_output),
    .io_passthrough(mac_2_27_io_passthrough)
  );
  MAC mac_2_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_28_clock),
    .reset(mac_2_28_reset),
    .io_load(mac_2_28_io_load),
    .io_mulInput(mac_2_28_io_mulInput),
    .io_addInput(mac_2_28_io_addInput),
    .io_output(mac_2_28_io_output),
    .io_passthrough(mac_2_28_io_passthrough)
  );
  MAC mac_2_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_29_clock),
    .reset(mac_2_29_reset),
    .io_load(mac_2_29_io_load),
    .io_mulInput(mac_2_29_io_mulInput),
    .io_addInput(mac_2_29_io_addInput),
    .io_output(mac_2_29_io_output),
    .io_passthrough(mac_2_29_io_passthrough)
  );
  MAC mac_2_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_30_clock),
    .reset(mac_2_30_reset),
    .io_load(mac_2_30_io_load),
    .io_mulInput(mac_2_30_io_mulInput),
    .io_addInput(mac_2_30_io_addInput),
    .io_output(mac_2_30_io_output),
    .io_passthrough(mac_2_30_io_passthrough)
  );
  MAC mac_2_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_2_31_clock),
    .reset(mac_2_31_reset),
    .io_load(mac_2_31_io_load),
    .io_mulInput(mac_2_31_io_mulInput),
    .io_addInput(mac_2_31_io_addInput),
    .io_output(mac_2_31_io_output),
    .io_passthrough(mac_2_31_io_passthrough)
  );
  MAC mac_3_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_0_clock),
    .reset(mac_3_0_reset),
    .io_load(mac_3_0_io_load),
    .io_mulInput(mac_3_0_io_mulInput),
    .io_addInput(mac_3_0_io_addInput),
    .io_output(mac_3_0_io_output),
    .io_passthrough(mac_3_0_io_passthrough)
  );
  MAC mac_3_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_1_clock),
    .reset(mac_3_1_reset),
    .io_load(mac_3_1_io_load),
    .io_mulInput(mac_3_1_io_mulInput),
    .io_addInput(mac_3_1_io_addInput),
    .io_output(mac_3_1_io_output),
    .io_passthrough(mac_3_1_io_passthrough)
  );
  MAC mac_3_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_2_clock),
    .reset(mac_3_2_reset),
    .io_load(mac_3_2_io_load),
    .io_mulInput(mac_3_2_io_mulInput),
    .io_addInput(mac_3_2_io_addInput),
    .io_output(mac_3_2_io_output),
    .io_passthrough(mac_3_2_io_passthrough)
  );
  MAC mac_3_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_3_clock),
    .reset(mac_3_3_reset),
    .io_load(mac_3_3_io_load),
    .io_mulInput(mac_3_3_io_mulInput),
    .io_addInput(mac_3_3_io_addInput),
    .io_output(mac_3_3_io_output),
    .io_passthrough(mac_3_3_io_passthrough)
  );
  MAC mac_3_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_4_clock),
    .reset(mac_3_4_reset),
    .io_load(mac_3_4_io_load),
    .io_mulInput(mac_3_4_io_mulInput),
    .io_addInput(mac_3_4_io_addInput),
    .io_output(mac_3_4_io_output),
    .io_passthrough(mac_3_4_io_passthrough)
  );
  MAC mac_3_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_5_clock),
    .reset(mac_3_5_reset),
    .io_load(mac_3_5_io_load),
    .io_mulInput(mac_3_5_io_mulInput),
    .io_addInput(mac_3_5_io_addInput),
    .io_output(mac_3_5_io_output),
    .io_passthrough(mac_3_5_io_passthrough)
  );
  MAC mac_3_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_6_clock),
    .reset(mac_3_6_reset),
    .io_load(mac_3_6_io_load),
    .io_mulInput(mac_3_6_io_mulInput),
    .io_addInput(mac_3_6_io_addInput),
    .io_output(mac_3_6_io_output),
    .io_passthrough(mac_3_6_io_passthrough)
  );
  MAC mac_3_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_7_clock),
    .reset(mac_3_7_reset),
    .io_load(mac_3_7_io_load),
    .io_mulInput(mac_3_7_io_mulInput),
    .io_addInput(mac_3_7_io_addInput),
    .io_output(mac_3_7_io_output),
    .io_passthrough(mac_3_7_io_passthrough)
  );
  MAC mac_3_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_8_clock),
    .reset(mac_3_8_reset),
    .io_load(mac_3_8_io_load),
    .io_mulInput(mac_3_8_io_mulInput),
    .io_addInput(mac_3_8_io_addInput),
    .io_output(mac_3_8_io_output),
    .io_passthrough(mac_3_8_io_passthrough)
  );
  MAC mac_3_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_9_clock),
    .reset(mac_3_9_reset),
    .io_load(mac_3_9_io_load),
    .io_mulInput(mac_3_9_io_mulInput),
    .io_addInput(mac_3_9_io_addInput),
    .io_output(mac_3_9_io_output),
    .io_passthrough(mac_3_9_io_passthrough)
  );
  MAC mac_3_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_10_clock),
    .reset(mac_3_10_reset),
    .io_load(mac_3_10_io_load),
    .io_mulInput(mac_3_10_io_mulInput),
    .io_addInput(mac_3_10_io_addInput),
    .io_output(mac_3_10_io_output),
    .io_passthrough(mac_3_10_io_passthrough)
  );
  MAC mac_3_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_11_clock),
    .reset(mac_3_11_reset),
    .io_load(mac_3_11_io_load),
    .io_mulInput(mac_3_11_io_mulInput),
    .io_addInput(mac_3_11_io_addInput),
    .io_output(mac_3_11_io_output),
    .io_passthrough(mac_3_11_io_passthrough)
  );
  MAC mac_3_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_12_clock),
    .reset(mac_3_12_reset),
    .io_load(mac_3_12_io_load),
    .io_mulInput(mac_3_12_io_mulInput),
    .io_addInput(mac_3_12_io_addInput),
    .io_output(mac_3_12_io_output),
    .io_passthrough(mac_3_12_io_passthrough)
  );
  MAC mac_3_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_13_clock),
    .reset(mac_3_13_reset),
    .io_load(mac_3_13_io_load),
    .io_mulInput(mac_3_13_io_mulInput),
    .io_addInput(mac_3_13_io_addInput),
    .io_output(mac_3_13_io_output),
    .io_passthrough(mac_3_13_io_passthrough)
  );
  MAC mac_3_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_14_clock),
    .reset(mac_3_14_reset),
    .io_load(mac_3_14_io_load),
    .io_mulInput(mac_3_14_io_mulInput),
    .io_addInput(mac_3_14_io_addInput),
    .io_output(mac_3_14_io_output),
    .io_passthrough(mac_3_14_io_passthrough)
  );
  MAC mac_3_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_15_clock),
    .reset(mac_3_15_reset),
    .io_load(mac_3_15_io_load),
    .io_mulInput(mac_3_15_io_mulInput),
    .io_addInput(mac_3_15_io_addInput),
    .io_output(mac_3_15_io_output),
    .io_passthrough(mac_3_15_io_passthrough)
  );
  MAC mac_3_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_16_clock),
    .reset(mac_3_16_reset),
    .io_load(mac_3_16_io_load),
    .io_mulInput(mac_3_16_io_mulInput),
    .io_addInput(mac_3_16_io_addInput),
    .io_output(mac_3_16_io_output),
    .io_passthrough(mac_3_16_io_passthrough)
  );
  MAC mac_3_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_17_clock),
    .reset(mac_3_17_reset),
    .io_load(mac_3_17_io_load),
    .io_mulInput(mac_3_17_io_mulInput),
    .io_addInput(mac_3_17_io_addInput),
    .io_output(mac_3_17_io_output),
    .io_passthrough(mac_3_17_io_passthrough)
  );
  MAC mac_3_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_18_clock),
    .reset(mac_3_18_reset),
    .io_load(mac_3_18_io_load),
    .io_mulInput(mac_3_18_io_mulInput),
    .io_addInput(mac_3_18_io_addInput),
    .io_output(mac_3_18_io_output),
    .io_passthrough(mac_3_18_io_passthrough)
  );
  MAC mac_3_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_19_clock),
    .reset(mac_3_19_reset),
    .io_load(mac_3_19_io_load),
    .io_mulInput(mac_3_19_io_mulInput),
    .io_addInput(mac_3_19_io_addInput),
    .io_output(mac_3_19_io_output),
    .io_passthrough(mac_3_19_io_passthrough)
  );
  MAC mac_3_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_20_clock),
    .reset(mac_3_20_reset),
    .io_load(mac_3_20_io_load),
    .io_mulInput(mac_3_20_io_mulInput),
    .io_addInput(mac_3_20_io_addInput),
    .io_output(mac_3_20_io_output),
    .io_passthrough(mac_3_20_io_passthrough)
  );
  MAC mac_3_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_21_clock),
    .reset(mac_3_21_reset),
    .io_load(mac_3_21_io_load),
    .io_mulInput(mac_3_21_io_mulInput),
    .io_addInput(mac_3_21_io_addInput),
    .io_output(mac_3_21_io_output),
    .io_passthrough(mac_3_21_io_passthrough)
  );
  MAC mac_3_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_22_clock),
    .reset(mac_3_22_reset),
    .io_load(mac_3_22_io_load),
    .io_mulInput(mac_3_22_io_mulInput),
    .io_addInput(mac_3_22_io_addInput),
    .io_output(mac_3_22_io_output),
    .io_passthrough(mac_3_22_io_passthrough)
  );
  MAC mac_3_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_23_clock),
    .reset(mac_3_23_reset),
    .io_load(mac_3_23_io_load),
    .io_mulInput(mac_3_23_io_mulInput),
    .io_addInput(mac_3_23_io_addInput),
    .io_output(mac_3_23_io_output),
    .io_passthrough(mac_3_23_io_passthrough)
  );
  MAC mac_3_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_24_clock),
    .reset(mac_3_24_reset),
    .io_load(mac_3_24_io_load),
    .io_mulInput(mac_3_24_io_mulInput),
    .io_addInput(mac_3_24_io_addInput),
    .io_output(mac_3_24_io_output),
    .io_passthrough(mac_3_24_io_passthrough)
  );
  MAC mac_3_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_25_clock),
    .reset(mac_3_25_reset),
    .io_load(mac_3_25_io_load),
    .io_mulInput(mac_3_25_io_mulInput),
    .io_addInput(mac_3_25_io_addInput),
    .io_output(mac_3_25_io_output),
    .io_passthrough(mac_3_25_io_passthrough)
  );
  MAC mac_3_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_26_clock),
    .reset(mac_3_26_reset),
    .io_load(mac_3_26_io_load),
    .io_mulInput(mac_3_26_io_mulInput),
    .io_addInput(mac_3_26_io_addInput),
    .io_output(mac_3_26_io_output),
    .io_passthrough(mac_3_26_io_passthrough)
  );
  MAC mac_3_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_27_clock),
    .reset(mac_3_27_reset),
    .io_load(mac_3_27_io_load),
    .io_mulInput(mac_3_27_io_mulInput),
    .io_addInput(mac_3_27_io_addInput),
    .io_output(mac_3_27_io_output),
    .io_passthrough(mac_3_27_io_passthrough)
  );
  MAC mac_3_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_28_clock),
    .reset(mac_3_28_reset),
    .io_load(mac_3_28_io_load),
    .io_mulInput(mac_3_28_io_mulInput),
    .io_addInput(mac_3_28_io_addInput),
    .io_output(mac_3_28_io_output),
    .io_passthrough(mac_3_28_io_passthrough)
  );
  MAC mac_3_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_29_clock),
    .reset(mac_3_29_reset),
    .io_load(mac_3_29_io_load),
    .io_mulInput(mac_3_29_io_mulInput),
    .io_addInput(mac_3_29_io_addInput),
    .io_output(mac_3_29_io_output),
    .io_passthrough(mac_3_29_io_passthrough)
  );
  MAC mac_3_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_30_clock),
    .reset(mac_3_30_reset),
    .io_load(mac_3_30_io_load),
    .io_mulInput(mac_3_30_io_mulInput),
    .io_addInput(mac_3_30_io_addInput),
    .io_output(mac_3_30_io_output),
    .io_passthrough(mac_3_30_io_passthrough)
  );
  MAC mac_3_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_3_31_clock),
    .reset(mac_3_31_reset),
    .io_load(mac_3_31_io_load),
    .io_mulInput(mac_3_31_io_mulInput),
    .io_addInput(mac_3_31_io_addInput),
    .io_output(mac_3_31_io_output),
    .io_passthrough(mac_3_31_io_passthrough)
  );
  MAC mac_4_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_0_clock),
    .reset(mac_4_0_reset),
    .io_load(mac_4_0_io_load),
    .io_mulInput(mac_4_0_io_mulInput),
    .io_addInput(mac_4_0_io_addInput),
    .io_output(mac_4_0_io_output),
    .io_passthrough(mac_4_0_io_passthrough)
  );
  MAC mac_4_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_1_clock),
    .reset(mac_4_1_reset),
    .io_load(mac_4_1_io_load),
    .io_mulInput(mac_4_1_io_mulInput),
    .io_addInput(mac_4_1_io_addInput),
    .io_output(mac_4_1_io_output),
    .io_passthrough(mac_4_1_io_passthrough)
  );
  MAC mac_4_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_2_clock),
    .reset(mac_4_2_reset),
    .io_load(mac_4_2_io_load),
    .io_mulInput(mac_4_2_io_mulInput),
    .io_addInput(mac_4_2_io_addInput),
    .io_output(mac_4_2_io_output),
    .io_passthrough(mac_4_2_io_passthrough)
  );
  MAC mac_4_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_3_clock),
    .reset(mac_4_3_reset),
    .io_load(mac_4_3_io_load),
    .io_mulInput(mac_4_3_io_mulInput),
    .io_addInput(mac_4_3_io_addInput),
    .io_output(mac_4_3_io_output),
    .io_passthrough(mac_4_3_io_passthrough)
  );
  MAC mac_4_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_4_clock),
    .reset(mac_4_4_reset),
    .io_load(mac_4_4_io_load),
    .io_mulInput(mac_4_4_io_mulInput),
    .io_addInput(mac_4_4_io_addInput),
    .io_output(mac_4_4_io_output),
    .io_passthrough(mac_4_4_io_passthrough)
  );
  MAC mac_4_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_5_clock),
    .reset(mac_4_5_reset),
    .io_load(mac_4_5_io_load),
    .io_mulInput(mac_4_5_io_mulInput),
    .io_addInput(mac_4_5_io_addInput),
    .io_output(mac_4_5_io_output),
    .io_passthrough(mac_4_5_io_passthrough)
  );
  MAC mac_4_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_6_clock),
    .reset(mac_4_6_reset),
    .io_load(mac_4_6_io_load),
    .io_mulInput(mac_4_6_io_mulInput),
    .io_addInput(mac_4_6_io_addInput),
    .io_output(mac_4_6_io_output),
    .io_passthrough(mac_4_6_io_passthrough)
  );
  MAC mac_4_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_7_clock),
    .reset(mac_4_7_reset),
    .io_load(mac_4_7_io_load),
    .io_mulInput(mac_4_7_io_mulInput),
    .io_addInput(mac_4_7_io_addInput),
    .io_output(mac_4_7_io_output),
    .io_passthrough(mac_4_7_io_passthrough)
  );
  MAC mac_4_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_8_clock),
    .reset(mac_4_8_reset),
    .io_load(mac_4_8_io_load),
    .io_mulInput(mac_4_8_io_mulInput),
    .io_addInput(mac_4_8_io_addInput),
    .io_output(mac_4_8_io_output),
    .io_passthrough(mac_4_8_io_passthrough)
  );
  MAC mac_4_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_9_clock),
    .reset(mac_4_9_reset),
    .io_load(mac_4_9_io_load),
    .io_mulInput(mac_4_9_io_mulInput),
    .io_addInput(mac_4_9_io_addInput),
    .io_output(mac_4_9_io_output),
    .io_passthrough(mac_4_9_io_passthrough)
  );
  MAC mac_4_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_10_clock),
    .reset(mac_4_10_reset),
    .io_load(mac_4_10_io_load),
    .io_mulInput(mac_4_10_io_mulInput),
    .io_addInput(mac_4_10_io_addInput),
    .io_output(mac_4_10_io_output),
    .io_passthrough(mac_4_10_io_passthrough)
  );
  MAC mac_4_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_11_clock),
    .reset(mac_4_11_reset),
    .io_load(mac_4_11_io_load),
    .io_mulInput(mac_4_11_io_mulInput),
    .io_addInput(mac_4_11_io_addInput),
    .io_output(mac_4_11_io_output),
    .io_passthrough(mac_4_11_io_passthrough)
  );
  MAC mac_4_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_12_clock),
    .reset(mac_4_12_reset),
    .io_load(mac_4_12_io_load),
    .io_mulInput(mac_4_12_io_mulInput),
    .io_addInput(mac_4_12_io_addInput),
    .io_output(mac_4_12_io_output),
    .io_passthrough(mac_4_12_io_passthrough)
  );
  MAC mac_4_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_13_clock),
    .reset(mac_4_13_reset),
    .io_load(mac_4_13_io_load),
    .io_mulInput(mac_4_13_io_mulInput),
    .io_addInput(mac_4_13_io_addInput),
    .io_output(mac_4_13_io_output),
    .io_passthrough(mac_4_13_io_passthrough)
  );
  MAC mac_4_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_14_clock),
    .reset(mac_4_14_reset),
    .io_load(mac_4_14_io_load),
    .io_mulInput(mac_4_14_io_mulInput),
    .io_addInput(mac_4_14_io_addInput),
    .io_output(mac_4_14_io_output),
    .io_passthrough(mac_4_14_io_passthrough)
  );
  MAC mac_4_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_15_clock),
    .reset(mac_4_15_reset),
    .io_load(mac_4_15_io_load),
    .io_mulInput(mac_4_15_io_mulInput),
    .io_addInput(mac_4_15_io_addInput),
    .io_output(mac_4_15_io_output),
    .io_passthrough(mac_4_15_io_passthrough)
  );
  MAC mac_4_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_16_clock),
    .reset(mac_4_16_reset),
    .io_load(mac_4_16_io_load),
    .io_mulInput(mac_4_16_io_mulInput),
    .io_addInput(mac_4_16_io_addInput),
    .io_output(mac_4_16_io_output),
    .io_passthrough(mac_4_16_io_passthrough)
  );
  MAC mac_4_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_17_clock),
    .reset(mac_4_17_reset),
    .io_load(mac_4_17_io_load),
    .io_mulInput(mac_4_17_io_mulInput),
    .io_addInput(mac_4_17_io_addInput),
    .io_output(mac_4_17_io_output),
    .io_passthrough(mac_4_17_io_passthrough)
  );
  MAC mac_4_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_18_clock),
    .reset(mac_4_18_reset),
    .io_load(mac_4_18_io_load),
    .io_mulInput(mac_4_18_io_mulInput),
    .io_addInput(mac_4_18_io_addInput),
    .io_output(mac_4_18_io_output),
    .io_passthrough(mac_4_18_io_passthrough)
  );
  MAC mac_4_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_19_clock),
    .reset(mac_4_19_reset),
    .io_load(mac_4_19_io_load),
    .io_mulInput(mac_4_19_io_mulInput),
    .io_addInput(mac_4_19_io_addInput),
    .io_output(mac_4_19_io_output),
    .io_passthrough(mac_4_19_io_passthrough)
  );
  MAC mac_4_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_20_clock),
    .reset(mac_4_20_reset),
    .io_load(mac_4_20_io_load),
    .io_mulInput(mac_4_20_io_mulInput),
    .io_addInput(mac_4_20_io_addInput),
    .io_output(mac_4_20_io_output),
    .io_passthrough(mac_4_20_io_passthrough)
  );
  MAC mac_4_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_21_clock),
    .reset(mac_4_21_reset),
    .io_load(mac_4_21_io_load),
    .io_mulInput(mac_4_21_io_mulInput),
    .io_addInput(mac_4_21_io_addInput),
    .io_output(mac_4_21_io_output),
    .io_passthrough(mac_4_21_io_passthrough)
  );
  MAC mac_4_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_22_clock),
    .reset(mac_4_22_reset),
    .io_load(mac_4_22_io_load),
    .io_mulInput(mac_4_22_io_mulInput),
    .io_addInput(mac_4_22_io_addInput),
    .io_output(mac_4_22_io_output),
    .io_passthrough(mac_4_22_io_passthrough)
  );
  MAC mac_4_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_23_clock),
    .reset(mac_4_23_reset),
    .io_load(mac_4_23_io_load),
    .io_mulInput(mac_4_23_io_mulInput),
    .io_addInput(mac_4_23_io_addInput),
    .io_output(mac_4_23_io_output),
    .io_passthrough(mac_4_23_io_passthrough)
  );
  MAC mac_4_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_24_clock),
    .reset(mac_4_24_reset),
    .io_load(mac_4_24_io_load),
    .io_mulInput(mac_4_24_io_mulInput),
    .io_addInput(mac_4_24_io_addInput),
    .io_output(mac_4_24_io_output),
    .io_passthrough(mac_4_24_io_passthrough)
  );
  MAC mac_4_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_25_clock),
    .reset(mac_4_25_reset),
    .io_load(mac_4_25_io_load),
    .io_mulInput(mac_4_25_io_mulInput),
    .io_addInput(mac_4_25_io_addInput),
    .io_output(mac_4_25_io_output),
    .io_passthrough(mac_4_25_io_passthrough)
  );
  MAC mac_4_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_26_clock),
    .reset(mac_4_26_reset),
    .io_load(mac_4_26_io_load),
    .io_mulInput(mac_4_26_io_mulInput),
    .io_addInput(mac_4_26_io_addInput),
    .io_output(mac_4_26_io_output),
    .io_passthrough(mac_4_26_io_passthrough)
  );
  MAC mac_4_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_27_clock),
    .reset(mac_4_27_reset),
    .io_load(mac_4_27_io_load),
    .io_mulInput(mac_4_27_io_mulInput),
    .io_addInput(mac_4_27_io_addInput),
    .io_output(mac_4_27_io_output),
    .io_passthrough(mac_4_27_io_passthrough)
  );
  MAC mac_4_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_28_clock),
    .reset(mac_4_28_reset),
    .io_load(mac_4_28_io_load),
    .io_mulInput(mac_4_28_io_mulInput),
    .io_addInput(mac_4_28_io_addInput),
    .io_output(mac_4_28_io_output),
    .io_passthrough(mac_4_28_io_passthrough)
  );
  MAC mac_4_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_29_clock),
    .reset(mac_4_29_reset),
    .io_load(mac_4_29_io_load),
    .io_mulInput(mac_4_29_io_mulInput),
    .io_addInput(mac_4_29_io_addInput),
    .io_output(mac_4_29_io_output),
    .io_passthrough(mac_4_29_io_passthrough)
  );
  MAC mac_4_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_30_clock),
    .reset(mac_4_30_reset),
    .io_load(mac_4_30_io_load),
    .io_mulInput(mac_4_30_io_mulInput),
    .io_addInput(mac_4_30_io_addInput),
    .io_output(mac_4_30_io_output),
    .io_passthrough(mac_4_30_io_passthrough)
  );
  MAC mac_4_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_4_31_clock),
    .reset(mac_4_31_reset),
    .io_load(mac_4_31_io_load),
    .io_mulInput(mac_4_31_io_mulInput),
    .io_addInput(mac_4_31_io_addInput),
    .io_output(mac_4_31_io_output),
    .io_passthrough(mac_4_31_io_passthrough)
  );
  MAC mac_5_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_0_clock),
    .reset(mac_5_0_reset),
    .io_load(mac_5_0_io_load),
    .io_mulInput(mac_5_0_io_mulInput),
    .io_addInput(mac_5_0_io_addInput),
    .io_output(mac_5_0_io_output),
    .io_passthrough(mac_5_0_io_passthrough)
  );
  MAC mac_5_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_1_clock),
    .reset(mac_5_1_reset),
    .io_load(mac_5_1_io_load),
    .io_mulInput(mac_5_1_io_mulInput),
    .io_addInput(mac_5_1_io_addInput),
    .io_output(mac_5_1_io_output),
    .io_passthrough(mac_5_1_io_passthrough)
  );
  MAC mac_5_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_2_clock),
    .reset(mac_5_2_reset),
    .io_load(mac_5_2_io_load),
    .io_mulInput(mac_5_2_io_mulInput),
    .io_addInput(mac_5_2_io_addInput),
    .io_output(mac_5_2_io_output),
    .io_passthrough(mac_5_2_io_passthrough)
  );
  MAC mac_5_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_3_clock),
    .reset(mac_5_3_reset),
    .io_load(mac_5_3_io_load),
    .io_mulInput(mac_5_3_io_mulInput),
    .io_addInput(mac_5_3_io_addInput),
    .io_output(mac_5_3_io_output),
    .io_passthrough(mac_5_3_io_passthrough)
  );
  MAC mac_5_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_4_clock),
    .reset(mac_5_4_reset),
    .io_load(mac_5_4_io_load),
    .io_mulInput(mac_5_4_io_mulInput),
    .io_addInput(mac_5_4_io_addInput),
    .io_output(mac_5_4_io_output),
    .io_passthrough(mac_5_4_io_passthrough)
  );
  MAC mac_5_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_5_clock),
    .reset(mac_5_5_reset),
    .io_load(mac_5_5_io_load),
    .io_mulInput(mac_5_5_io_mulInput),
    .io_addInput(mac_5_5_io_addInput),
    .io_output(mac_5_5_io_output),
    .io_passthrough(mac_5_5_io_passthrough)
  );
  MAC mac_5_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_6_clock),
    .reset(mac_5_6_reset),
    .io_load(mac_5_6_io_load),
    .io_mulInput(mac_5_6_io_mulInput),
    .io_addInput(mac_5_6_io_addInput),
    .io_output(mac_5_6_io_output),
    .io_passthrough(mac_5_6_io_passthrough)
  );
  MAC mac_5_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_7_clock),
    .reset(mac_5_7_reset),
    .io_load(mac_5_7_io_load),
    .io_mulInput(mac_5_7_io_mulInput),
    .io_addInput(mac_5_7_io_addInput),
    .io_output(mac_5_7_io_output),
    .io_passthrough(mac_5_7_io_passthrough)
  );
  MAC mac_5_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_8_clock),
    .reset(mac_5_8_reset),
    .io_load(mac_5_8_io_load),
    .io_mulInput(mac_5_8_io_mulInput),
    .io_addInput(mac_5_8_io_addInput),
    .io_output(mac_5_8_io_output),
    .io_passthrough(mac_5_8_io_passthrough)
  );
  MAC mac_5_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_9_clock),
    .reset(mac_5_9_reset),
    .io_load(mac_5_9_io_load),
    .io_mulInput(mac_5_9_io_mulInput),
    .io_addInput(mac_5_9_io_addInput),
    .io_output(mac_5_9_io_output),
    .io_passthrough(mac_5_9_io_passthrough)
  );
  MAC mac_5_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_10_clock),
    .reset(mac_5_10_reset),
    .io_load(mac_5_10_io_load),
    .io_mulInput(mac_5_10_io_mulInput),
    .io_addInput(mac_5_10_io_addInput),
    .io_output(mac_5_10_io_output),
    .io_passthrough(mac_5_10_io_passthrough)
  );
  MAC mac_5_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_11_clock),
    .reset(mac_5_11_reset),
    .io_load(mac_5_11_io_load),
    .io_mulInput(mac_5_11_io_mulInput),
    .io_addInput(mac_5_11_io_addInput),
    .io_output(mac_5_11_io_output),
    .io_passthrough(mac_5_11_io_passthrough)
  );
  MAC mac_5_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_12_clock),
    .reset(mac_5_12_reset),
    .io_load(mac_5_12_io_load),
    .io_mulInput(mac_5_12_io_mulInput),
    .io_addInput(mac_5_12_io_addInput),
    .io_output(mac_5_12_io_output),
    .io_passthrough(mac_5_12_io_passthrough)
  );
  MAC mac_5_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_13_clock),
    .reset(mac_5_13_reset),
    .io_load(mac_5_13_io_load),
    .io_mulInput(mac_5_13_io_mulInput),
    .io_addInput(mac_5_13_io_addInput),
    .io_output(mac_5_13_io_output),
    .io_passthrough(mac_5_13_io_passthrough)
  );
  MAC mac_5_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_14_clock),
    .reset(mac_5_14_reset),
    .io_load(mac_5_14_io_load),
    .io_mulInput(mac_5_14_io_mulInput),
    .io_addInput(mac_5_14_io_addInput),
    .io_output(mac_5_14_io_output),
    .io_passthrough(mac_5_14_io_passthrough)
  );
  MAC mac_5_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_15_clock),
    .reset(mac_5_15_reset),
    .io_load(mac_5_15_io_load),
    .io_mulInput(mac_5_15_io_mulInput),
    .io_addInput(mac_5_15_io_addInput),
    .io_output(mac_5_15_io_output),
    .io_passthrough(mac_5_15_io_passthrough)
  );
  MAC mac_5_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_16_clock),
    .reset(mac_5_16_reset),
    .io_load(mac_5_16_io_load),
    .io_mulInput(mac_5_16_io_mulInput),
    .io_addInput(mac_5_16_io_addInput),
    .io_output(mac_5_16_io_output),
    .io_passthrough(mac_5_16_io_passthrough)
  );
  MAC mac_5_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_17_clock),
    .reset(mac_5_17_reset),
    .io_load(mac_5_17_io_load),
    .io_mulInput(mac_5_17_io_mulInput),
    .io_addInput(mac_5_17_io_addInput),
    .io_output(mac_5_17_io_output),
    .io_passthrough(mac_5_17_io_passthrough)
  );
  MAC mac_5_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_18_clock),
    .reset(mac_5_18_reset),
    .io_load(mac_5_18_io_load),
    .io_mulInput(mac_5_18_io_mulInput),
    .io_addInput(mac_5_18_io_addInput),
    .io_output(mac_5_18_io_output),
    .io_passthrough(mac_5_18_io_passthrough)
  );
  MAC mac_5_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_19_clock),
    .reset(mac_5_19_reset),
    .io_load(mac_5_19_io_load),
    .io_mulInput(mac_5_19_io_mulInput),
    .io_addInput(mac_5_19_io_addInput),
    .io_output(mac_5_19_io_output),
    .io_passthrough(mac_5_19_io_passthrough)
  );
  MAC mac_5_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_20_clock),
    .reset(mac_5_20_reset),
    .io_load(mac_5_20_io_load),
    .io_mulInput(mac_5_20_io_mulInput),
    .io_addInput(mac_5_20_io_addInput),
    .io_output(mac_5_20_io_output),
    .io_passthrough(mac_5_20_io_passthrough)
  );
  MAC mac_5_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_21_clock),
    .reset(mac_5_21_reset),
    .io_load(mac_5_21_io_load),
    .io_mulInput(mac_5_21_io_mulInput),
    .io_addInput(mac_5_21_io_addInput),
    .io_output(mac_5_21_io_output),
    .io_passthrough(mac_5_21_io_passthrough)
  );
  MAC mac_5_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_22_clock),
    .reset(mac_5_22_reset),
    .io_load(mac_5_22_io_load),
    .io_mulInput(mac_5_22_io_mulInput),
    .io_addInput(mac_5_22_io_addInput),
    .io_output(mac_5_22_io_output),
    .io_passthrough(mac_5_22_io_passthrough)
  );
  MAC mac_5_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_23_clock),
    .reset(mac_5_23_reset),
    .io_load(mac_5_23_io_load),
    .io_mulInput(mac_5_23_io_mulInput),
    .io_addInput(mac_5_23_io_addInput),
    .io_output(mac_5_23_io_output),
    .io_passthrough(mac_5_23_io_passthrough)
  );
  MAC mac_5_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_24_clock),
    .reset(mac_5_24_reset),
    .io_load(mac_5_24_io_load),
    .io_mulInput(mac_5_24_io_mulInput),
    .io_addInput(mac_5_24_io_addInput),
    .io_output(mac_5_24_io_output),
    .io_passthrough(mac_5_24_io_passthrough)
  );
  MAC mac_5_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_25_clock),
    .reset(mac_5_25_reset),
    .io_load(mac_5_25_io_load),
    .io_mulInput(mac_5_25_io_mulInput),
    .io_addInput(mac_5_25_io_addInput),
    .io_output(mac_5_25_io_output),
    .io_passthrough(mac_5_25_io_passthrough)
  );
  MAC mac_5_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_26_clock),
    .reset(mac_5_26_reset),
    .io_load(mac_5_26_io_load),
    .io_mulInput(mac_5_26_io_mulInput),
    .io_addInput(mac_5_26_io_addInput),
    .io_output(mac_5_26_io_output),
    .io_passthrough(mac_5_26_io_passthrough)
  );
  MAC mac_5_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_27_clock),
    .reset(mac_5_27_reset),
    .io_load(mac_5_27_io_load),
    .io_mulInput(mac_5_27_io_mulInput),
    .io_addInput(mac_5_27_io_addInput),
    .io_output(mac_5_27_io_output),
    .io_passthrough(mac_5_27_io_passthrough)
  );
  MAC mac_5_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_28_clock),
    .reset(mac_5_28_reset),
    .io_load(mac_5_28_io_load),
    .io_mulInput(mac_5_28_io_mulInput),
    .io_addInput(mac_5_28_io_addInput),
    .io_output(mac_5_28_io_output),
    .io_passthrough(mac_5_28_io_passthrough)
  );
  MAC mac_5_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_29_clock),
    .reset(mac_5_29_reset),
    .io_load(mac_5_29_io_load),
    .io_mulInput(mac_5_29_io_mulInput),
    .io_addInput(mac_5_29_io_addInput),
    .io_output(mac_5_29_io_output),
    .io_passthrough(mac_5_29_io_passthrough)
  );
  MAC mac_5_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_30_clock),
    .reset(mac_5_30_reset),
    .io_load(mac_5_30_io_load),
    .io_mulInput(mac_5_30_io_mulInput),
    .io_addInput(mac_5_30_io_addInput),
    .io_output(mac_5_30_io_output),
    .io_passthrough(mac_5_30_io_passthrough)
  );
  MAC mac_5_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_5_31_clock),
    .reset(mac_5_31_reset),
    .io_load(mac_5_31_io_load),
    .io_mulInput(mac_5_31_io_mulInput),
    .io_addInput(mac_5_31_io_addInput),
    .io_output(mac_5_31_io_output),
    .io_passthrough(mac_5_31_io_passthrough)
  );
  MAC mac_6_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_0_clock),
    .reset(mac_6_0_reset),
    .io_load(mac_6_0_io_load),
    .io_mulInput(mac_6_0_io_mulInput),
    .io_addInput(mac_6_0_io_addInput),
    .io_output(mac_6_0_io_output),
    .io_passthrough(mac_6_0_io_passthrough)
  );
  MAC mac_6_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_1_clock),
    .reset(mac_6_1_reset),
    .io_load(mac_6_1_io_load),
    .io_mulInput(mac_6_1_io_mulInput),
    .io_addInput(mac_6_1_io_addInput),
    .io_output(mac_6_1_io_output),
    .io_passthrough(mac_6_1_io_passthrough)
  );
  MAC mac_6_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_2_clock),
    .reset(mac_6_2_reset),
    .io_load(mac_6_2_io_load),
    .io_mulInput(mac_6_2_io_mulInput),
    .io_addInput(mac_6_2_io_addInput),
    .io_output(mac_6_2_io_output),
    .io_passthrough(mac_6_2_io_passthrough)
  );
  MAC mac_6_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_3_clock),
    .reset(mac_6_3_reset),
    .io_load(mac_6_3_io_load),
    .io_mulInput(mac_6_3_io_mulInput),
    .io_addInput(mac_6_3_io_addInput),
    .io_output(mac_6_3_io_output),
    .io_passthrough(mac_6_3_io_passthrough)
  );
  MAC mac_6_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_4_clock),
    .reset(mac_6_4_reset),
    .io_load(mac_6_4_io_load),
    .io_mulInput(mac_6_4_io_mulInput),
    .io_addInput(mac_6_4_io_addInput),
    .io_output(mac_6_4_io_output),
    .io_passthrough(mac_6_4_io_passthrough)
  );
  MAC mac_6_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_5_clock),
    .reset(mac_6_5_reset),
    .io_load(mac_6_5_io_load),
    .io_mulInput(mac_6_5_io_mulInput),
    .io_addInput(mac_6_5_io_addInput),
    .io_output(mac_6_5_io_output),
    .io_passthrough(mac_6_5_io_passthrough)
  );
  MAC mac_6_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_6_clock),
    .reset(mac_6_6_reset),
    .io_load(mac_6_6_io_load),
    .io_mulInput(mac_6_6_io_mulInput),
    .io_addInput(mac_6_6_io_addInput),
    .io_output(mac_6_6_io_output),
    .io_passthrough(mac_6_6_io_passthrough)
  );
  MAC mac_6_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_7_clock),
    .reset(mac_6_7_reset),
    .io_load(mac_6_7_io_load),
    .io_mulInput(mac_6_7_io_mulInput),
    .io_addInput(mac_6_7_io_addInput),
    .io_output(mac_6_7_io_output),
    .io_passthrough(mac_6_7_io_passthrough)
  );
  MAC mac_6_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_8_clock),
    .reset(mac_6_8_reset),
    .io_load(mac_6_8_io_load),
    .io_mulInput(mac_6_8_io_mulInput),
    .io_addInput(mac_6_8_io_addInput),
    .io_output(mac_6_8_io_output),
    .io_passthrough(mac_6_8_io_passthrough)
  );
  MAC mac_6_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_9_clock),
    .reset(mac_6_9_reset),
    .io_load(mac_6_9_io_load),
    .io_mulInput(mac_6_9_io_mulInput),
    .io_addInput(mac_6_9_io_addInput),
    .io_output(mac_6_9_io_output),
    .io_passthrough(mac_6_9_io_passthrough)
  );
  MAC mac_6_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_10_clock),
    .reset(mac_6_10_reset),
    .io_load(mac_6_10_io_load),
    .io_mulInput(mac_6_10_io_mulInput),
    .io_addInput(mac_6_10_io_addInput),
    .io_output(mac_6_10_io_output),
    .io_passthrough(mac_6_10_io_passthrough)
  );
  MAC mac_6_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_11_clock),
    .reset(mac_6_11_reset),
    .io_load(mac_6_11_io_load),
    .io_mulInput(mac_6_11_io_mulInput),
    .io_addInput(mac_6_11_io_addInput),
    .io_output(mac_6_11_io_output),
    .io_passthrough(mac_6_11_io_passthrough)
  );
  MAC mac_6_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_12_clock),
    .reset(mac_6_12_reset),
    .io_load(mac_6_12_io_load),
    .io_mulInput(mac_6_12_io_mulInput),
    .io_addInput(mac_6_12_io_addInput),
    .io_output(mac_6_12_io_output),
    .io_passthrough(mac_6_12_io_passthrough)
  );
  MAC mac_6_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_13_clock),
    .reset(mac_6_13_reset),
    .io_load(mac_6_13_io_load),
    .io_mulInput(mac_6_13_io_mulInput),
    .io_addInput(mac_6_13_io_addInput),
    .io_output(mac_6_13_io_output),
    .io_passthrough(mac_6_13_io_passthrough)
  );
  MAC mac_6_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_14_clock),
    .reset(mac_6_14_reset),
    .io_load(mac_6_14_io_load),
    .io_mulInput(mac_6_14_io_mulInput),
    .io_addInput(mac_6_14_io_addInput),
    .io_output(mac_6_14_io_output),
    .io_passthrough(mac_6_14_io_passthrough)
  );
  MAC mac_6_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_15_clock),
    .reset(mac_6_15_reset),
    .io_load(mac_6_15_io_load),
    .io_mulInput(mac_6_15_io_mulInput),
    .io_addInput(mac_6_15_io_addInput),
    .io_output(mac_6_15_io_output),
    .io_passthrough(mac_6_15_io_passthrough)
  );
  MAC mac_6_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_16_clock),
    .reset(mac_6_16_reset),
    .io_load(mac_6_16_io_load),
    .io_mulInput(mac_6_16_io_mulInput),
    .io_addInput(mac_6_16_io_addInput),
    .io_output(mac_6_16_io_output),
    .io_passthrough(mac_6_16_io_passthrough)
  );
  MAC mac_6_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_17_clock),
    .reset(mac_6_17_reset),
    .io_load(mac_6_17_io_load),
    .io_mulInput(mac_6_17_io_mulInput),
    .io_addInput(mac_6_17_io_addInput),
    .io_output(mac_6_17_io_output),
    .io_passthrough(mac_6_17_io_passthrough)
  );
  MAC mac_6_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_18_clock),
    .reset(mac_6_18_reset),
    .io_load(mac_6_18_io_load),
    .io_mulInput(mac_6_18_io_mulInput),
    .io_addInput(mac_6_18_io_addInput),
    .io_output(mac_6_18_io_output),
    .io_passthrough(mac_6_18_io_passthrough)
  );
  MAC mac_6_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_19_clock),
    .reset(mac_6_19_reset),
    .io_load(mac_6_19_io_load),
    .io_mulInput(mac_6_19_io_mulInput),
    .io_addInput(mac_6_19_io_addInput),
    .io_output(mac_6_19_io_output),
    .io_passthrough(mac_6_19_io_passthrough)
  );
  MAC mac_6_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_20_clock),
    .reset(mac_6_20_reset),
    .io_load(mac_6_20_io_load),
    .io_mulInput(mac_6_20_io_mulInput),
    .io_addInput(mac_6_20_io_addInput),
    .io_output(mac_6_20_io_output),
    .io_passthrough(mac_6_20_io_passthrough)
  );
  MAC mac_6_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_21_clock),
    .reset(mac_6_21_reset),
    .io_load(mac_6_21_io_load),
    .io_mulInput(mac_6_21_io_mulInput),
    .io_addInput(mac_6_21_io_addInput),
    .io_output(mac_6_21_io_output),
    .io_passthrough(mac_6_21_io_passthrough)
  );
  MAC mac_6_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_22_clock),
    .reset(mac_6_22_reset),
    .io_load(mac_6_22_io_load),
    .io_mulInput(mac_6_22_io_mulInput),
    .io_addInput(mac_6_22_io_addInput),
    .io_output(mac_6_22_io_output),
    .io_passthrough(mac_6_22_io_passthrough)
  );
  MAC mac_6_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_23_clock),
    .reset(mac_6_23_reset),
    .io_load(mac_6_23_io_load),
    .io_mulInput(mac_6_23_io_mulInput),
    .io_addInput(mac_6_23_io_addInput),
    .io_output(mac_6_23_io_output),
    .io_passthrough(mac_6_23_io_passthrough)
  );
  MAC mac_6_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_24_clock),
    .reset(mac_6_24_reset),
    .io_load(mac_6_24_io_load),
    .io_mulInput(mac_6_24_io_mulInput),
    .io_addInput(mac_6_24_io_addInput),
    .io_output(mac_6_24_io_output),
    .io_passthrough(mac_6_24_io_passthrough)
  );
  MAC mac_6_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_25_clock),
    .reset(mac_6_25_reset),
    .io_load(mac_6_25_io_load),
    .io_mulInput(mac_6_25_io_mulInput),
    .io_addInput(mac_6_25_io_addInput),
    .io_output(mac_6_25_io_output),
    .io_passthrough(mac_6_25_io_passthrough)
  );
  MAC mac_6_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_26_clock),
    .reset(mac_6_26_reset),
    .io_load(mac_6_26_io_load),
    .io_mulInput(mac_6_26_io_mulInput),
    .io_addInput(mac_6_26_io_addInput),
    .io_output(mac_6_26_io_output),
    .io_passthrough(mac_6_26_io_passthrough)
  );
  MAC mac_6_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_27_clock),
    .reset(mac_6_27_reset),
    .io_load(mac_6_27_io_load),
    .io_mulInput(mac_6_27_io_mulInput),
    .io_addInput(mac_6_27_io_addInput),
    .io_output(mac_6_27_io_output),
    .io_passthrough(mac_6_27_io_passthrough)
  );
  MAC mac_6_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_28_clock),
    .reset(mac_6_28_reset),
    .io_load(mac_6_28_io_load),
    .io_mulInput(mac_6_28_io_mulInput),
    .io_addInput(mac_6_28_io_addInput),
    .io_output(mac_6_28_io_output),
    .io_passthrough(mac_6_28_io_passthrough)
  );
  MAC mac_6_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_29_clock),
    .reset(mac_6_29_reset),
    .io_load(mac_6_29_io_load),
    .io_mulInput(mac_6_29_io_mulInput),
    .io_addInput(mac_6_29_io_addInput),
    .io_output(mac_6_29_io_output),
    .io_passthrough(mac_6_29_io_passthrough)
  );
  MAC mac_6_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_30_clock),
    .reset(mac_6_30_reset),
    .io_load(mac_6_30_io_load),
    .io_mulInput(mac_6_30_io_mulInput),
    .io_addInput(mac_6_30_io_addInput),
    .io_output(mac_6_30_io_output),
    .io_passthrough(mac_6_30_io_passthrough)
  );
  MAC mac_6_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_6_31_clock),
    .reset(mac_6_31_reset),
    .io_load(mac_6_31_io_load),
    .io_mulInput(mac_6_31_io_mulInput),
    .io_addInput(mac_6_31_io_addInput),
    .io_output(mac_6_31_io_output),
    .io_passthrough(mac_6_31_io_passthrough)
  );
  MAC mac_7_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_0_clock),
    .reset(mac_7_0_reset),
    .io_load(mac_7_0_io_load),
    .io_mulInput(mac_7_0_io_mulInput),
    .io_addInput(mac_7_0_io_addInput),
    .io_output(mac_7_0_io_output),
    .io_passthrough(mac_7_0_io_passthrough)
  );
  MAC mac_7_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_1_clock),
    .reset(mac_7_1_reset),
    .io_load(mac_7_1_io_load),
    .io_mulInput(mac_7_1_io_mulInput),
    .io_addInput(mac_7_1_io_addInput),
    .io_output(mac_7_1_io_output),
    .io_passthrough(mac_7_1_io_passthrough)
  );
  MAC mac_7_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_2_clock),
    .reset(mac_7_2_reset),
    .io_load(mac_7_2_io_load),
    .io_mulInput(mac_7_2_io_mulInput),
    .io_addInput(mac_7_2_io_addInput),
    .io_output(mac_7_2_io_output),
    .io_passthrough(mac_7_2_io_passthrough)
  );
  MAC mac_7_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_3_clock),
    .reset(mac_7_3_reset),
    .io_load(mac_7_3_io_load),
    .io_mulInput(mac_7_3_io_mulInput),
    .io_addInput(mac_7_3_io_addInput),
    .io_output(mac_7_3_io_output),
    .io_passthrough(mac_7_3_io_passthrough)
  );
  MAC mac_7_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_4_clock),
    .reset(mac_7_4_reset),
    .io_load(mac_7_4_io_load),
    .io_mulInput(mac_7_4_io_mulInput),
    .io_addInput(mac_7_4_io_addInput),
    .io_output(mac_7_4_io_output),
    .io_passthrough(mac_7_4_io_passthrough)
  );
  MAC mac_7_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_5_clock),
    .reset(mac_7_5_reset),
    .io_load(mac_7_5_io_load),
    .io_mulInput(mac_7_5_io_mulInput),
    .io_addInput(mac_7_5_io_addInput),
    .io_output(mac_7_5_io_output),
    .io_passthrough(mac_7_5_io_passthrough)
  );
  MAC mac_7_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_6_clock),
    .reset(mac_7_6_reset),
    .io_load(mac_7_6_io_load),
    .io_mulInput(mac_7_6_io_mulInput),
    .io_addInput(mac_7_6_io_addInput),
    .io_output(mac_7_6_io_output),
    .io_passthrough(mac_7_6_io_passthrough)
  );
  MAC mac_7_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_7_clock),
    .reset(mac_7_7_reset),
    .io_load(mac_7_7_io_load),
    .io_mulInput(mac_7_7_io_mulInput),
    .io_addInput(mac_7_7_io_addInput),
    .io_output(mac_7_7_io_output),
    .io_passthrough(mac_7_7_io_passthrough)
  );
  MAC mac_7_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_8_clock),
    .reset(mac_7_8_reset),
    .io_load(mac_7_8_io_load),
    .io_mulInput(mac_7_8_io_mulInput),
    .io_addInput(mac_7_8_io_addInput),
    .io_output(mac_7_8_io_output),
    .io_passthrough(mac_7_8_io_passthrough)
  );
  MAC mac_7_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_9_clock),
    .reset(mac_7_9_reset),
    .io_load(mac_7_9_io_load),
    .io_mulInput(mac_7_9_io_mulInput),
    .io_addInput(mac_7_9_io_addInput),
    .io_output(mac_7_9_io_output),
    .io_passthrough(mac_7_9_io_passthrough)
  );
  MAC mac_7_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_10_clock),
    .reset(mac_7_10_reset),
    .io_load(mac_7_10_io_load),
    .io_mulInput(mac_7_10_io_mulInput),
    .io_addInput(mac_7_10_io_addInput),
    .io_output(mac_7_10_io_output),
    .io_passthrough(mac_7_10_io_passthrough)
  );
  MAC mac_7_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_11_clock),
    .reset(mac_7_11_reset),
    .io_load(mac_7_11_io_load),
    .io_mulInput(mac_7_11_io_mulInput),
    .io_addInput(mac_7_11_io_addInput),
    .io_output(mac_7_11_io_output),
    .io_passthrough(mac_7_11_io_passthrough)
  );
  MAC mac_7_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_12_clock),
    .reset(mac_7_12_reset),
    .io_load(mac_7_12_io_load),
    .io_mulInput(mac_7_12_io_mulInput),
    .io_addInput(mac_7_12_io_addInput),
    .io_output(mac_7_12_io_output),
    .io_passthrough(mac_7_12_io_passthrough)
  );
  MAC mac_7_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_13_clock),
    .reset(mac_7_13_reset),
    .io_load(mac_7_13_io_load),
    .io_mulInput(mac_7_13_io_mulInput),
    .io_addInput(mac_7_13_io_addInput),
    .io_output(mac_7_13_io_output),
    .io_passthrough(mac_7_13_io_passthrough)
  );
  MAC mac_7_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_14_clock),
    .reset(mac_7_14_reset),
    .io_load(mac_7_14_io_load),
    .io_mulInput(mac_7_14_io_mulInput),
    .io_addInput(mac_7_14_io_addInput),
    .io_output(mac_7_14_io_output),
    .io_passthrough(mac_7_14_io_passthrough)
  );
  MAC mac_7_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_15_clock),
    .reset(mac_7_15_reset),
    .io_load(mac_7_15_io_load),
    .io_mulInput(mac_7_15_io_mulInput),
    .io_addInput(mac_7_15_io_addInput),
    .io_output(mac_7_15_io_output),
    .io_passthrough(mac_7_15_io_passthrough)
  );
  MAC mac_7_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_16_clock),
    .reset(mac_7_16_reset),
    .io_load(mac_7_16_io_load),
    .io_mulInput(mac_7_16_io_mulInput),
    .io_addInput(mac_7_16_io_addInput),
    .io_output(mac_7_16_io_output),
    .io_passthrough(mac_7_16_io_passthrough)
  );
  MAC mac_7_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_17_clock),
    .reset(mac_7_17_reset),
    .io_load(mac_7_17_io_load),
    .io_mulInput(mac_7_17_io_mulInput),
    .io_addInput(mac_7_17_io_addInput),
    .io_output(mac_7_17_io_output),
    .io_passthrough(mac_7_17_io_passthrough)
  );
  MAC mac_7_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_18_clock),
    .reset(mac_7_18_reset),
    .io_load(mac_7_18_io_load),
    .io_mulInput(mac_7_18_io_mulInput),
    .io_addInput(mac_7_18_io_addInput),
    .io_output(mac_7_18_io_output),
    .io_passthrough(mac_7_18_io_passthrough)
  );
  MAC mac_7_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_19_clock),
    .reset(mac_7_19_reset),
    .io_load(mac_7_19_io_load),
    .io_mulInput(mac_7_19_io_mulInput),
    .io_addInput(mac_7_19_io_addInput),
    .io_output(mac_7_19_io_output),
    .io_passthrough(mac_7_19_io_passthrough)
  );
  MAC mac_7_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_20_clock),
    .reset(mac_7_20_reset),
    .io_load(mac_7_20_io_load),
    .io_mulInput(mac_7_20_io_mulInput),
    .io_addInput(mac_7_20_io_addInput),
    .io_output(mac_7_20_io_output),
    .io_passthrough(mac_7_20_io_passthrough)
  );
  MAC mac_7_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_21_clock),
    .reset(mac_7_21_reset),
    .io_load(mac_7_21_io_load),
    .io_mulInput(mac_7_21_io_mulInput),
    .io_addInput(mac_7_21_io_addInput),
    .io_output(mac_7_21_io_output),
    .io_passthrough(mac_7_21_io_passthrough)
  );
  MAC mac_7_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_22_clock),
    .reset(mac_7_22_reset),
    .io_load(mac_7_22_io_load),
    .io_mulInput(mac_7_22_io_mulInput),
    .io_addInput(mac_7_22_io_addInput),
    .io_output(mac_7_22_io_output),
    .io_passthrough(mac_7_22_io_passthrough)
  );
  MAC mac_7_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_23_clock),
    .reset(mac_7_23_reset),
    .io_load(mac_7_23_io_load),
    .io_mulInput(mac_7_23_io_mulInput),
    .io_addInput(mac_7_23_io_addInput),
    .io_output(mac_7_23_io_output),
    .io_passthrough(mac_7_23_io_passthrough)
  );
  MAC mac_7_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_24_clock),
    .reset(mac_7_24_reset),
    .io_load(mac_7_24_io_load),
    .io_mulInput(mac_7_24_io_mulInput),
    .io_addInput(mac_7_24_io_addInput),
    .io_output(mac_7_24_io_output),
    .io_passthrough(mac_7_24_io_passthrough)
  );
  MAC mac_7_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_25_clock),
    .reset(mac_7_25_reset),
    .io_load(mac_7_25_io_load),
    .io_mulInput(mac_7_25_io_mulInput),
    .io_addInput(mac_7_25_io_addInput),
    .io_output(mac_7_25_io_output),
    .io_passthrough(mac_7_25_io_passthrough)
  );
  MAC mac_7_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_26_clock),
    .reset(mac_7_26_reset),
    .io_load(mac_7_26_io_load),
    .io_mulInput(mac_7_26_io_mulInput),
    .io_addInput(mac_7_26_io_addInput),
    .io_output(mac_7_26_io_output),
    .io_passthrough(mac_7_26_io_passthrough)
  );
  MAC mac_7_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_27_clock),
    .reset(mac_7_27_reset),
    .io_load(mac_7_27_io_load),
    .io_mulInput(mac_7_27_io_mulInput),
    .io_addInput(mac_7_27_io_addInput),
    .io_output(mac_7_27_io_output),
    .io_passthrough(mac_7_27_io_passthrough)
  );
  MAC mac_7_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_28_clock),
    .reset(mac_7_28_reset),
    .io_load(mac_7_28_io_load),
    .io_mulInput(mac_7_28_io_mulInput),
    .io_addInput(mac_7_28_io_addInput),
    .io_output(mac_7_28_io_output),
    .io_passthrough(mac_7_28_io_passthrough)
  );
  MAC mac_7_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_29_clock),
    .reset(mac_7_29_reset),
    .io_load(mac_7_29_io_load),
    .io_mulInput(mac_7_29_io_mulInput),
    .io_addInput(mac_7_29_io_addInput),
    .io_output(mac_7_29_io_output),
    .io_passthrough(mac_7_29_io_passthrough)
  );
  MAC mac_7_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_30_clock),
    .reset(mac_7_30_reset),
    .io_load(mac_7_30_io_load),
    .io_mulInput(mac_7_30_io_mulInput),
    .io_addInput(mac_7_30_io_addInput),
    .io_output(mac_7_30_io_output),
    .io_passthrough(mac_7_30_io_passthrough)
  );
  MAC mac_7_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_7_31_clock),
    .reset(mac_7_31_reset),
    .io_load(mac_7_31_io_load),
    .io_mulInput(mac_7_31_io_mulInput),
    .io_addInput(mac_7_31_io_addInput),
    .io_output(mac_7_31_io_output),
    .io_passthrough(mac_7_31_io_passthrough)
  );
  MAC mac_8_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_0_clock),
    .reset(mac_8_0_reset),
    .io_load(mac_8_0_io_load),
    .io_mulInput(mac_8_0_io_mulInput),
    .io_addInput(mac_8_0_io_addInput),
    .io_output(mac_8_0_io_output),
    .io_passthrough(mac_8_0_io_passthrough)
  );
  MAC mac_8_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_1_clock),
    .reset(mac_8_1_reset),
    .io_load(mac_8_1_io_load),
    .io_mulInput(mac_8_1_io_mulInput),
    .io_addInput(mac_8_1_io_addInput),
    .io_output(mac_8_1_io_output),
    .io_passthrough(mac_8_1_io_passthrough)
  );
  MAC mac_8_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_2_clock),
    .reset(mac_8_2_reset),
    .io_load(mac_8_2_io_load),
    .io_mulInput(mac_8_2_io_mulInput),
    .io_addInput(mac_8_2_io_addInput),
    .io_output(mac_8_2_io_output),
    .io_passthrough(mac_8_2_io_passthrough)
  );
  MAC mac_8_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_3_clock),
    .reset(mac_8_3_reset),
    .io_load(mac_8_3_io_load),
    .io_mulInput(mac_8_3_io_mulInput),
    .io_addInput(mac_8_3_io_addInput),
    .io_output(mac_8_3_io_output),
    .io_passthrough(mac_8_3_io_passthrough)
  );
  MAC mac_8_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_4_clock),
    .reset(mac_8_4_reset),
    .io_load(mac_8_4_io_load),
    .io_mulInput(mac_8_4_io_mulInput),
    .io_addInput(mac_8_4_io_addInput),
    .io_output(mac_8_4_io_output),
    .io_passthrough(mac_8_4_io_passthrough)
  );
  MAC mac_8_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_5_clock),
    .reset(mac_8_5_reset),
    .io_load(mac_8_5_io_load),
    .io_mulInput(mac_8_5_io_mulInput),
    .io_addInput(mac_8_5_io_addInput),
    .io_output(mac_8_5_io_output),
    .io_passthrough(mac_8_5_io_passthrough)
  );
  MAC mac_8_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_6_clock),
    .reset(mac_8_6_reset),
    .io_load(mac_8_6_io_load),
    .io_mulInput(mac_8_6_io_mulInput),
    .io_addInput(mac_8_6_io_addInput),
    .io_output(mac_8_6_io_output),
    .io_passthrough(mac_8_6_io_passthrough)
  );
  MAC mac_8_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_7_clock),
    .reset(mac_8_7_reset),
    .io_load(mac_8_7_io_load),
    .io_mulInput(mac_8_7_io_mulInput),
    .io_addInput(mac_8_7_io_addInput),
    .io_output(mac_8_7_io_output),
    .io_passthrough(mac_8_7_io_passthrough)
  );
  MAC mac_8_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_8_clock),
    .reset(mac_8_8_reset),
    .io_load(mac_8_8_io_load),
    .io_mulInput(mac_8_8_io_mulInput),
    .io_addInput(mac_8_8_io_addInput),
    .io_output(mac_8_8_io_output),
    .io_passthrough(mac_8_8_io_passthrough)
  );
  MAC mac_8_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_9_clock),
    .reset(mac_8_9_reset),
    .io_load(mac_8_9_io_load),
    .io_mulInput(mac_8_9_io_mulInput),
    .io_addInput(mac_8_9_io_addInput),
    .io_output(mac_8_9_io_output),
    .io_passthrough(mac_8_9_io_passthrough)
  );
  MAC mac_8_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_10_clock),
    .reset(mac_8_10_reset),
    .io_load(mac_8_10_io_load),
    .io_mulInput(mac_8_10_io_mulInput),
    .io_addInput(mac_8_10_io_addInput),
    .io_output(mac_8_10_io_output),
    .io_passthrough(mac_8_10_io_passthrough)
  );
  MAC mac_8_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_11_clock),
    .reset(mac_8_11_reset),
    .io_load(mac_8_11_io_load),
    .io_mulInput(mac_8_11_io_mulInput),
    .io_addInput(mac_8_11_io_addInput),
    .io_output(mac_8_11_io_output),
    .io_passthrough(mac_8_11_io_passthrough)
  );
  MAC mac_8_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_12_clock),
    .reset(mac_8_12_reset),
    .io_load(mac_8_12_io_load),
    .io_mulInput(mac_8_12_io_mulInput),
    .io_addInput(mac_8_12_io_addInput),
    .io_output(mac_8_12_io_output),
    .io_passthrough(mac_8_12_io_passthrough)
  );
  MAC mac_8_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_13_clock),
    .reset(mac_8_13_reset),
    .io_load(mac_8_13_io_load),
    .io_mulInput(mac_8_13_io_mulInput),
    .io_addInput(mac_8_13_io_addInput),
    .io_output(mac_8_13_io_output),
    .io_passthrough(mac_8_13_io_passthrough)
  );
  MAC mac_8_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_14_clock),
    .reset(mac_8_14_reset),
    .io_load(mac_8_14_io_load),
    .io_mulInput(mac_8_14_io_mulInput),
    .io_addInput(mac_8_14_io_addInput),
    .io_output(mac_8_14_io_output),
    .io_passthrough(mac_8_14_io_passthrough)
  );
  MAC mac_8_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_15_clock),
    .reset(mac_8_15_reset),
    .io_load(mac_8_15_io_load),
    .io_mulInput(mac_8_15_io_mulInput),
    .io_addInput(mac_8_15_io_addInput),
    .io_output(mac_8_15_io_output),
    .io_passthrough(mac_8_15_io_passthrough)
  );
  MAC mac_8_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_16_clock),
    .reset(mac_8_16_reset),
    .io_load(mac_8_16_io_load),
    .io_mulInput(mac_8_16_io_mulInput),
    .io_addInput(mac_8_16_io_addInput),
    .io_output(mac_8_16_io_output),
    .io_passthrough(mac_8_16_io_passthrough)
  );
  MAC mac_8_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_17_clock),
    .reset(mac_8_17_reset),
    .io_load(mac_8_17_io_load),
    .io_mulInput(mac_8_17_io_mulInput),
    .io_addInput(mac_8_17_io_addInput),
    .io_output(mac_8_17_io_output),
    .io_passthrough(mac_8_17_io_passthrough)
  );
  MAC mac_8_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_18_clock),
    .reset(mac_8_18_reset),
    .io_load(mac_8_18_io_load),
    .io_mulInput(mac_8_18_io_mulInput),
    .io_addInput(mac_8_18_io_addInput),
    .io_output(mac_8_18_io_output),
    .io_passthrough(mac_8_18_io_passthrough)
  );
  MAC mac_8_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_19_clock),
    .reset(mac_8_19_reset),
    .io_load(mac_8_19_io_load),
    .io_mulInput(mac_8_19_io_mulInput),
    .io_addInput(mac_8_19_io_addInput),
    .io_output(mac_8_19_io_output),
    .io_passthrough(mac_8_19_io_passthrough)
  );
  MAC mac_8_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_20_clock),
    .reset(mac_8_20_reset),
    .io_load(mac_8_20_io_load),
    .io_mulInput(mac_8_20_io_mulInput),
    .io_addInput(mac_8_20_io_addInput),
    .io_output(mac_8_20_io_output),
    .io_passthrough(mac_8_20_io_passthrough)
  );
  MAC mac_8_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_21_clock),
    .reset(mac_8_21_reset),
    .io_load(mac_8_21_io_load),
    .io_mulInput(mac_8_21_io_mulInput),
    .io_addInput(mac_8_21_io_addInput),
    .io_output(mac_8_21_io_output),
    .io_passthrough(mac_8_21_io_passthrough)
  );
  MAC mac_8_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_22_clock),
    .reset(mac_8_22_reset),
    .io_load(mac_8_22_io_load),
    .io_mulInput(mac_8_22_io_mulInput),
    .io_addInput(mac_8_22_io_addInput),
    .io_output(mac_8_22_io_output),
    .io_passthrough(mac_8_22_io_passthrough)
  );
  MAC mac_8_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_23_clock),
    .reset(mac_8_23_reset),
    .io_load(mac_8_23_io_load),
    .io_mulInput(mac_8_23_io_mulInput),
    .io_addInput(mac_8_23_io_addInput),
    .io_output(mac_8_23_io_output),
    .io_passthrough(mac_8_23_io_passthrough)
  );
  MAC mac_8_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_24_clock),
    .reset(mac_8_24_reset),
    .io_load(mac_8_24_io_load),
    .io_mulInput(mac_8_24_io_mulInput),
    .io_addInput(mac_8_24_io_addInput),
    .io_output(mac_8_24_io_output),
    .io_passthrough(mac_8_24_io_passthrough)
  );
  MAC mac_8_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_25_clock),
    .reset(mac_8_25_reset),
    .io_load(mac_8_25_io_load),
    .io_mulInput(mac_8_25_io_mulInput),
    .io_addInput(mac_8_25_io_addInput),
    .io_output(mac_8_25_io_output),
    .io_passthrough(mac_8_25_io_passthrough)
  );
  MAC mac_8_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_26_clock),
    .reset(mac_8_26_reset),
    .io_load(mac_8_26_io_load),
    .io_mulInput(mac_8_26_io_mulInput),
    .io_addInput(mac_8_26_io_addInput),
    .io_output(mac_8_26_io_output),
    .io_passthrough(mac_8_26_io_passthrough)
  );
  MAC mac_8_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_27_clock),
    .reset(mac_8_27_reset),
    .io_load(mac_8_27_io_load),
    .io_mulInput(mac_8_27_io_mulInput),
    .io_addInput(mac_8_27_io_addInput),
    .io_output(mac_8_27_io_output),
    .io_passthrough(mac_8_27_io_passthrough)
  );
  MAC mac_8_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_28_clock),
    .reset(mac_8_28_reset),
    .io_load(mac_8_28_io_load),
    .io_mulInput(mac_8_28_io_mulInput),
    .io_addInput(mac_8_28_io_addInput),
    .io_output(mac_8_28_io_output),
    .io_passthrough(mac_8_28_io_passthrough)
  );
  MAC mac_8_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_29_clock),
    .reset(mac_8_29_reset),
    .io_load(mac_8_29_io_load),
    .io_mulInput(mac_8_29_io_mulInput),
    .io_addInput(mac_8_29_io_addInput),
    .io_output(mac_8_29_io_output),
    .io_passthrough(mac_8_29_io_passthrough)
  );
  MAC mac_8_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_30_clock),
    .reset(mac_8_30_reset),
    .io_load(mac_8_30_io_load),
    .io_mulInput(mac_8_30_io_mulInput),
    .io_addInput(mac_8_30_io_addInput),
    .io_output(mac_8_30_io_output),
    .io_passthrough(mac_8_30_io_passthrough)
  );
  MAC mac_8_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_8_31_clock),
    .reset(mac_8_31_reset),
    .io_load(mac_8_31_io_load),
    .io_mulInput(mac_8_31_io_mulInput),
    .io_addInput(mac_8_31_io_addInput),
    .io_output(mac_8_31_io_output),
    .io_passthrough(mac_8_31_io_passthrough)
  );
  MAC mac_9_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_0_clock),
    .reset(mac_9_0_reset),
    .io_load(mac_9_0_io_load),
    .io_mulInput(mac_9_0_io_mulInput),
    .io_addInput(mac_9_0_io_addInput),
    .io_output(mac_9_0_io_output),
    .io_passthrough(mac_9_0_io_passthrough)
  );
  MAC mac_9_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_1_clock),
    .reset(mac_9_1_reset),
    .io_load(mac_9_1_io_load),
    .io_mulInput(mac_9_1_io_mulInput),
    .io_addInput(mac_9_1_io_addInput),
    .io_output(mac_9_1_io_output),
    .io_passthrough(mac_9_1_io_passthrough)
  );
  MAC mac_9_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_2_clock),
    .reset(mac_9_2_reset),
    .io_load(mac_9_2_io_load),
    .io_mulInput(mac_9_2_io_mulInput),
    .io_addInput(mac_9_2_io_addInput),
    .io_output(mac_9_2_io_output),
    .io_passthrough(mac_9_2_io_passthrough)
  );
  MAC mac_9_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_3_clock),
    .reset(mac_9_3_reset),
    .io_load(mac_9_3_io_load),
    .io_mulInput(mac_9_3_io_mulInput),
    .io_addInput(mac_9_3_io_addInput),
    .io_output(mac_9_3_io_output),
    .io_passthrough(mac_9_3_io_passthrough)
  );
  MAC mac_9_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_4_clock),
    .reset(mac_9_4_reset),
    .io_load(mac_9_4_io_load),
    .io_mulInput(mac_9_4_io_mulInput),
    .io_addInput(mac_9_4_io_addInput),
    .io_output(mac_9_4_io_output),
    .io_passthrough(mac_9_4_io_passthrough)
  );
  MAC mac_9_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_5_clock),
    .reset(mac_9_5_reset),
    .io_load(mac_9_5_io_load),
    .io_mulInput(mac_9_5_io_mulInput),
    .io_addInput(mac_9_5_io_addInput),
    .io_output(mac_9_5_io_output),
    .io_passthrough(mac_9_5_io_passthrough)
  );
  MAC mac_9_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_6_clock),
    .reset(mac_9_6_reset),
    .io_load(mac_9_6_io_load),
    .io_mulInput(mac_9_6_io_mulInput),
    .io_addInput(mac_9_6_io_addInput),
    .io_output(mac_9_6_io_output),
    .io_passthrough(mac_9_6_io_passthrough)
  );
  MAC mac_9_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_7_clock),
    .reset(mac_9_7_reset),
    .io_load(mac_9_7_io_load),
    .io_mulInput(mac_9_7_io_mulInput),
    .io_addInput(mac_9_7_io_addInput),
    .io_output(mac_9_7_io_output),
    .io_passthrough(mac_9_7_io_passthrough)
  );
  MAC mac_9_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_8_clock),
    .reset(mac_9_8_reset),
    .io_load(mac_9_8_io_load),
    .io_mulInput(mac_9_8_io_mulInput),
    .io_addInput(mac_9_8_io_addInput),
    .io_output(mac_9_8_io_output),
    .io_passthrough(mac_9_8_io_passthrough)
  );
  MAC mac_9_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_9_clock),
    .reset(mac_9_9_reset),
    .io_load(mac_9_9_io_load),
    .io_mulInput(mac_9_9_io_mulInput),
    .io_addInput(mac_9_9_io_addInput),
    .io_output(mac_9_9_io_output),
    .io_passthrough(mac_9_9_io_passthrough)
  );
  MAC mac_9_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_10_clock),
    .reset(mac_9_10_reset),
    .io_load(mac_9_10_io_load),
    .io_mulInput(mac_9_10_io_mulInput),
    .io_addInput(mac_9_10_io_addInput),
    .io_output(mac_9_10_io_output),
    .io_passthrough(mac_9_10_io_passthrough)
  );
  MAC mac_9_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_11_clock),
    .reset(mac_9_11_reset),
    .io_load(mac_9_11_io_load),
    .io_mulInput(mac_9_11_io_mulInput),
    .io_addInput(mac_9_11_io_addInput),
    .io_output(mac_9_11_io_output),
    .io_passthrough(mac_9_11_io_passthrough)
  );
  MAC mac_9_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_12_clock),
    .reset(mac_9_12_reset),
    .io_load(mac_9_12_io_load),
    .io_mulInput(mac_9_12_io_mulInput),
    .io_addInput(mac_9_12_io_addInput),
    .io_output(mac_9_12_io_output),
    .io_passthrough(mac_9_12_io_passthrough)
  );
  MAC mac_9_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_13_clock),
    .reset(mac_9_13_reset),
    .io_load(mac_9_13_io_load),
    .io_mulInput(mac_9_13_io_mulInput),
    .io_addInput(mac_9_13_io_addInput),
    .io_output(mac_9_13_io_output),
    .io_passthrough(mac_9_13_io_passthrough)
  );
  MAC mac_9_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_14_clock),
    .reset(mac_9_14_reset),
    .io_load(mac_9_14_io_load),
    .io_mulInput(mac_9_14_io_mulInput),
    .io_addInput(mac_9_14_io_addInput),
    .io_output(mac_9_14_io_output),
    .io_passthrough(mac_9_14_io_passthrough)
  );
  MAC mac_9_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_15_clock),
    .reset(mac_9_15_reset),
    .io_load(mac_9_15_io_load),
    .io_mulInput(mac_9_15_io_mulInput),
    .io_addInput(mac_9_15_io_addInput),
    .io_output(mac_9_15_io_output),
    .io_passthrough(mac_9_15_io_passthrough)
  );
  MAC mac_9_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_16_clock),
    .reset(mac_9_16_reset),
    .io_load(mac_9_16_io_load),
    .io_mulInput(mac_9_16_io_mulInput),
    .io_addInput(mac_9_16_io_addInput),
    .io_output(mac_9_16_io_output),
    .io_passthrough(mac_9_16_io_passthrough)
  );
  MAC mac_9_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_17_clock),
    .reset(mac_9_17_reset),
    .io_load(mac_9_17_io_load),
    .io_mulInput(mac_9_17_io_mulInput),
    .io_addInput(mac_9_17_io_addInput),
    .io_output(mac_9_17_io_output),
    .io_passthrough(mac_9_17_io_passthrough)
  );
  MAC mac_9_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_18_clock),
    .reset(mac_9_18_reset),
    .io_load(mac_9_18_io_load),
    .io_mulInput(mac_9_18_io_mulInput),
    .io_addInput(mac_9_18_io_addInput),
    .io_output(mac_9_18_io_output),
    .io_passthrough(mac_9_18_io_passthrough)
  );
  MAC mac_9_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_19_clock),
    .reset(mac_9_19_reset),
    .io_load(mac_9_19_io_load),
    .io_mulInput(mac_9_19_io_mulInput),
    .io_addInput(mac_9_19_io_addInput),
    .io_output(mac_9_19_io_output),
    .io_passthrough(mac_9_19_io_passthrough)
  );
  MAC mac_9_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_20_clock),
    .reset(mac_9_20_reset),
    .io_load(mac_9_20_io_load),
    .io_mulInput(mac_9_20_io_mulInput),
    .io_addInput(mac_9_20_io_addInput),
    .io_output(mac_9_20_io_output),
    .io_passthrough(mac_9_20_io_passthrough)
  );
  MAC mac_9_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_21_clock),
    .reset(mac_9_21_reset),
    .io_load(mac_9_21_io_load),
    .io_mulInput(mac_9_21_io_mulInput),
    .io_addInput(mac_9_21_io_addInput),
    .io_output(mac_9_21_io_output),
    .io_passthrough(mac_9_21_io_passthrough)
  );
  MAC mac_9_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_22_clock),
    .reset(mac_9_22_reset),
    .io_load(mac_9_22_io_load),
    .io_mulInput(mac_9_22_io_mulInput),
    .io_addInput(mac_9_22_io_addInput),
    .io_output(mac_9_22_io_output),
    .io_passthrough(mac_9_22_io_passthrough)
  );
  MAC mac_9_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_23_clock),
    .reset(mac_9_23_reset),
    .io_load(mac_9_23_io_load),
    .io_mulInput(mac_9_23_io_mulInput),
    .io_addInput(mac_9_23_io_addInput),
    .io_output(mac_9_23_io_output),
    .io_passthrough(mac_9_23_io_passthrough)
  );
  MAC mac_9_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_24_clock),
    .reset(mac_9_24_reset),
    .io_load(mac_9_24_io_load),
    .io_mulInput(mac_9_24_io_mulInput),
    .io_addInput(mac_9_24_io_addInput),
    .io_output(mac_9_24_io_output),
    .io_passthrough(mac_9_24_io_passthrough)
  );
  MAC mac_9_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_25_clock),
    .reset(mac_9_25_reset),
    .io_load(mac_9_25_io_load),
    .io_mulInput(mac_9_25_io_mulInput),
    .io_addInput(mac_9_25_io_addInput),
    .io_output(mac_9_25_io_output),
    .io_passthrough(mac_9_25_io_passthrough)
  );
  MAC mac_9_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_26_clock),
    .reset(mac_9_26_reset),
    .io_load(mac_9_26_io_load),
    .io_mulInput(mac_9_26_io_mulInput),
    .io_addInput(mac_9_26_io_addInput),
    .io_output(mac_9_26_io_output),
    .io_passthrough(mac_9_26_io_passthrough)
  );
  MAC mac_9_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_27_clock),
    .reset(mac_9_27_reset),
    .io_load(mac_9_27_io_load),
    .io_mulInput(mac_9_27_io_mulInput),
    .io_addInput(mac_9_27_io_addInput),
    .io_output(mac_9_27_io_output),
    .io_passthrough(mac_9_27_io_passthrough)
  );
  MAC mac_9_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_28_clock),
    .reset(mac_9_28_reset),
    .io_load(mac_9_28_io_load),
    .io_mulInput(mac_9_28_io_mulInput),
    .io_addInput(mac_9_28_io_addInput),
    .io_output(mac_9_28_io_output),
    .io_passthrough(mac_9_28_io_passthrough)
  );
  MAC mac_9_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_29_clock),
    .reset(mac_9_29_reset),
    .io_load(mac_9_29_io_load),
    .io_mulInput(mac_9_29_io_mulInput),
    .io_addInput(mac_9_29_io_addInput),
    .io_output(mac_9_29_io_output),
    .io_passthrough(mac_9_29_io_passthrough)
  );
  MAC mac_9_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_30_clock),
    .reset(mac_9_30_reset),
    .io_load(mac_9_30_io_load),
    .io_mulInput(mac_9_30_io_mulInput),
    .io_addInput(mac_9_30_io_addInput),
    .io_output(mac_9_30_io_output),
    .io_passthrough(mac_9_30_io_passthrough)
  );
  MAC mac_9_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_9_31_clock),
    .reset(mac_9_31_reset),
    .io_load(mac_9_31_io_load),
    .io_mulInput(mac_9_31_io_mulInput),
    .io_addInput(mac_9_31_io_addInput),
    .io_output(mac_9_31_io_output),
    .io_passthrough(mac_9_31_io_passthrough)
  );
  MAC mac_10_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_0_clock),
    .reset(mac_10_0_reset),
    .io_load(mac_10_0_io_load),
    .io_mulInput(mac_10_0_io_mulInput),
    .io_addInput(mac_10_0_io_addInput),
    .io_output(mac_10_0_io_output),
    .io_passthrough(mac_10_0_io_passthrough)
  );
  MAC mac_10_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_1_clock),
    .reset(mac_10_1_reset),
    .io_load(mac_10_1_io_load),
    .io_mulInput(mac_10_1_io_mulInput),
    .io_addInput(mac_10_1_io_addInput),
    .io_output(mac_10_1_io_output),
    .io_passthrough(mac_10_1_io_passthrough)
  );
  MAC mac_10_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_2_clock),
    .reset(mac_10_2_reset),
    .io_load(mac_10_2_io_load),
    .io_mulInput(mac_10_2_io_mulInput),
    .io_addInput(mac_10_2_io_addInput),
    .io_output(mac_10_2_io_output),
    .io_passthrough(mac_10_2_io_passthrough)
  );
  MAC mac_10_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_3_clock),
    .reset(mac_10_3_reset),
    .io_load(mac_10_3_io_load),
    .io_mulInput(mac_10_3_io_mulInput),
    .io_addInput(mac_10_3_io_addInput),
    .io_output(mac_10_3_io_output),
    .io_passthrough(mac_10_3_io_passthrough)
  );
  MAC mac_10_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_4_clock),
    .reset(mac_10_4_reset),
    .io_load(mac_10_4_io_load),
    .io_mulInput(mac_10_4_io_mulInput),
    .io_addInput(mac_10_4_io_addInput),
    .io_output(mac_10_4_io_output),
    .io_passthrough(mac_10_4_io_passthrough)
  );
  MAC mac_10_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_5_clock),
    .reset(mac_10_5_reset),
    .io_load(mac_10_5_io_load),
    .io_mulInput(mac_10_5_io_mulInput),
    .io_addInput(mac_10_5_io_addInput),
    .io_output(mac_10_5_io_output),
    .io_passthrough(mac_10_5_io_passthrough)
  );
  MAC mac_10_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_6_clock),
    .reset(mac_10_6_reset),
    .io_load(mac_10_6_io_load),
    .io_mulInput(mac_10_6_io_mulInput),
    .io_addInput(mac_10_6_io_addInput),
    .io_output(mac_10_6_io_output),
    .io_passthrough(mac_10_6_io_passthrough)
  );
  MAC mac_10_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_7_clock),
    .reset(mac_10_7_reset),
    .io_load(mac_10_7_io_load),
    .io_mulInput(mac_10_7_io_mulInput),
    .io_addInput(mac_10_7_io_addInput),
    .io_output(mac_10_7_io_output),
    .io_passthrough(mac_10_7_io_passthrough)
  );
  MAC mac_10_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_8_clock),
    .reset(mac_10_8_reset),
    .io_load(mac_10_8_io_load),
    .io_mulInput(mac_10_8_io_mulInput),
    .io_addInput(mac_10_8_io_addInput),
    .io_output(mac_10_8_io_output),
    .io_passthrough(mac_10_8_io_passthrough)
  );
  MAC mac_10_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_9_clock),
    .reset(mac_10_9_reset),
    .io_load(mac_10_9_io_load),
    .io_mulInput(mac_10_9_io_mulInput),
    .io_addInput(mac_10_9_io_addInput),
    .io_output(mac_10_9_io_output),
    .io_passthrough(mac_10_9_io_passthrough)
  );
  MAC mac_10_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_10_clock),
    .reset(mac_10_10_reset),
    .io_load(mac_10_10_io_load),
    .io_mulInput(mac_10_10_io_mulInput),
    .io_addInput(mac_10_10_io_addInput),
    .io_output(mac_10_10_io_output),
    .io_passthrough(mac_10_10_io_passthrough)
  );
  MAC mac_10_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_11_clock),
    .reset(mac_10_11_reset),
    .io_load(mac_10_11_io_load),
    .io_mulInput(mac_10_11_io_mulInput),
    .io_addInput(mac_10_11_io_addInput),
    .io_output(mac_10_11_io_output),
    .io_passthrough(mac_10_11_io_passthrough)
  );
  MAC mac_10_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_12_clock),
    .reset(mac_10_12_reset),
    .io_load(mac_10_12_io_load),
    .io_mulInput(mac_10_12_io_mulInput),
    .io_addInput(mac_10_12_io_addInput),
    .io_output(mac_10_12_io_output),
    .io_passthrough(mac_10_12_io_passthrough)
  );
  MAC mac_10_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_13_clock),
    .reset(mac_10_13_reset),
    .io_load(mac_10_13_io_load),
    .io_mulInput(mac_10_13_io_mulInput),
    .io_addInput(mac_10_13_io_addInput),
    .io_output(mac_10_13_io_output),
    .io_passthrough(mac_10_13_io_passthrough)
  );
  MAC mac_10_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_14_clock),
    .reset(mac_10_14_reset),
    .io_load(mac_10_14_io_load),
    .io_mulInput(mac_10_14_io_mulInput),
    .io_addInput(mac_10_14_io_addInput),
    .io_output(mac_10_14_io_output),
    .io_passthrough(mac_10_14_io_passthrough)
  );
  MAC mac_10_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_15_clock),
    .reset(mac_10_15_reset),
    .io_load(mac_10_15_io_load),
    .io_mulInput(mac_10_15_io_mulInput),
    .io_addInput(mac_10_15_io_addInput),
    .io_output(mac_10_15_io_output),
    .io_passthrough(mac_10_15_io_passthrough)
  );
  MAC mac_10_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_16_clock),
    .reset(mac_10_16_reset),
    .io_load(mac_10_16_io_load),
    .io_mulInput(mac_10_16_io_mulInput),
    .io_addInput(mac_10_16_io_addInput),
    .io_output(mac_10_16_io_output),
    .io_passthrough(mac_10_16_io_passthrough)
  );
  MAC mac_10_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_17_clock),
    .reset(mac_10_17_reset),
    .io_load(mac_10_17_io_load),
    .io_mulInput(mac_10_17_io_mulInput),
    .io_addInput(mac_10_17_io_addInput),
    .io_output(mac_10_17_io_output),
    .io_passthrough(mac_10_17_io_passthrough)
  );
  MAC mac_10_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_18_clock),
    .reset(mac_10_18_reset),
    .io_load(mac_10_18_io_load),
    .io_mulInput(mac_10_18_io_mulInput),
    .io_addInput(mac_10_18_io_addInput),
    .io_output(mac_10_18_io_output),
    .io_passthrough(mac_10_18_io_passthrough)
  );
  MAC mac_10_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_19_clock),
    .reset(mac_10_19_reset),
    .io_load(mac_10_19_io_load),
    .io_mulInput(mac_10_19_io_mulInput),
    .io_addInput(mac_10_19_io_addInput),
    .io_output(mac_10_19_io_output),
    .io_passthrough(mac_10_19_io_passthrough)
  );
  MAC mac_10_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_20_clock),
    .reset(mac_10_20_reset),
    .io_load(mac_10_20_io_load),
    .io_mulInput(mac_10_20_io_mulInput),
    .io_addInput(mac_10_20_io_addInput),
    .io_output(mac_10_20_io_output),
    .io_passthrough(mac_10_20_io_passthrough)
  );
  MAC mac_10_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_21_clock),
    .reset(mac_10_21_reset),
    .io_load(mac_10_21_io_load),
    .io_mulInput(mac_10_21_io_mulInput),
    .io_addInput(mac_10_21_io_addInput),
    .io_output(mac_10_21_io_output),
    .io_passthrough(mac_10_21_io_passthrough)
  );
  MAC mac_10_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_22_clock),
    .reset(mac_10_22_reset),
    .io_load(mac_10_22_io_load),
    .io_mulInput(mac_10_22_io_mulInput),
    .io_addInput(mac_10_22_io_addInput),
    .io_output(mac_10_22_io_output),
    .io_passthrough(mac_10_22_io_passthrough)
  );
  MAC mac_10_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_23_clock),
    .reset(mac_10_23_reset),
    .io_load(mac_10_23_io_load),
    .io_mulInput(mac_10_23_io_mulInput),
    .io_addInput(mac_10_23_io_addInput),
    .io_output(mac_10_23_io_output),
    .io_passthrough(mac_10_23_io_passthrough)
  );
  MAC mac_10_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_24_clock),
    .reset(mac_10_24_reset),
    .io_load(mac_10_24_io_load),
    .io_mulInput(mac_10_24_io_mulInput),
    .io_addInput(mac_10_24_io_addInput),
    .io_output(mac_10_24_io_output),
    .io_passthrough(mac_10_24_io_passthrough)
  );
  MAC mac_10_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_25_clock),
    .reset(mac_10_25_reset),
    .io_load(mac_10_25_io_load),
    .io_mulInput(mac_10_25_io_mulInput),
    .io_addInput(mac_10_25_io_addInput),
    .io_output(mac_10_25_io_output),
    .io_passthrough(mac_10_25_io_passthrough)
  );
  MAC mac_10_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_26_clock),
    .reset(mac_10_26_reset),
    .io_load(mac_10_26_io_load),
    .io_mulInput(mac_10_26_io_mulInput),
    .io_addInput(mac_10_26_io_addInput),
    .io_output(mac_10_26_io_output),
    .io_passthrough(mac_10_26_io_passthrough)
  );
  MAC mac_10_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_27_clock),
    .reset(mac_10_27_reset),
    .io_load(mac_10_27_io_load),
    .io_mulInput(mac_10_27_io_mulInput),
    .io_addInput(mac_10_27_io_addInput),
    .io_output(mac_10_27_io_output),
    .io_passthrough(mac_10_27_io_passthrough)
  );
  MAC mac_10_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_28_clock),
    .reset(mac_10_28_reset),
    .io_load(mac_10_28_io_load),
    .io_mulInput(mac_10_28_io_mulInput),
    .io_addInput(mac_10_28_io_addInput),
    .io_output(mac_10_28_io_output),
    .io_passthrough(mac_10_28_io_passthrough)
  );
  MAC mac_10_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_29_clock),
    .reset(mac_10_29_reset),
    .io_load(mac_10_29_io_load),
    .io_mulInput(mac_10_29_io_mulInput),
    .io_addInput(mac_10_29_io_addInput),
    .io_output(mac_10_29_io_output),
    .io_passthrough(mac_10_29_io_passthrough)
  );
  MAC mac_10_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_30_clock),
    .reset(mac_10_30_reset),
    .io_load(mac_10_30_io_load),
    .io_mulInput(mac_10_30_io_mulInput),
    .io_addInput(mac_10_30_io_addInput),
    .io_output(mac_10_30_io_output),
    .io_passthrough(mac_10_30_io_passthrough)
  );
  MAC mac_10_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_10_31_clock),
    .reset(mac_10_31_reset),
    .io_load(mac_10_31_io_load),
    .io_mulInput(mac_10_31_io_mulInput),
    .io_addInput(mac_10_31_io_addInput),
    .io_output(mac_10_31_io_output),
    .io_passthrough(mac_10_31_io_passthrough)
  );
  MAC mac_11_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_0_clock),
    .reset(mac_11_0_reset),
    .io_load(mac_11_0_io_load),
    .io_mulInput(mac_11_0_io_mulInput),
    .io_addInput(mac_11_0_io_addInput),
    .io_output(mac_11_0_io_output),
    .io_passthrough(mac_11_0_io_passthrough)
  );
  MAC mac_11_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_1_clock),
    .reset(mac_11_1_reset),
    .io_load(mac_11_1_io_load),
    .io_mulInput(mac_11_1_io_mulInput),
    .io_addInput(mac_11_1_io_addInput),
    .io_output(mac_11_1_io_output),
    .io_passthrough(mac_11_1_io_passthrough)
  );
  MAC mac_11_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_2_clock),
    .reset(mac_11_2_reset),
    .io_load(mac_11_2_io_load),
    .io_mulInput(mac_11_2_io_mulInput),
    .io_addInput(mac_11_2_io_addInput),
    .io_output(mac_11_2_io_output),
    .io_passthrough(mac_11_2_io_passthrough)
  );
  MAC mac_11_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_3_clock),
    .reset(mac_11_3_reset),
    .io_load(mac_11_3_io_load),
    .io_mulInput(mac_11_3_io_mulInput),
    .io_addInput(mac_11_3_io_addInput),
    .io_output(mac_11_3_io_output),
    .io_passthrough(mac_11_3_io_passthrough)
  );
  MAC mac_11_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_4_clock),
    .reset(mac_11_4_reset),
    .io_load(mac_11_4_io_load),
    .io_mulInput(mac_11_4_io_mulInput),
    .io_addInput(mac_11_4_io_addInput),
    .io_output(mac_11_4_io_output),
    .io_passthrough(mac_11_4_io_passthrough)
  );
  MAC mac_11_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_5_clock),
    .reset(mac_11_5_reset),
    .io_load(mac_11_5_io_load),
    .io_mulInput(mac_11_5_io_mulInput),
    .io_addInput(mac_11_5_io_addInput),
    .io_output(mac_11_5_io_output),
    .io_passthrough(mac_11_5_io_passthrough)
  );
  MAC mac_11_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_6_clock),
    .reset(mac_11_6_reset),
    .io_load(mac_11_6_io_load),
    .io_mulInput(mac_11_6_io_mulInput),
    .io_addInput(mac_11_6_io_addInput),
    .io_output(mac_11_6_io_output),
    .io_passthrough(mac_11_6_io_passthrough)
  );
  MAC mac_11_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_7_clock),
    .reset(mac_11_7_reset),
    .io_load(mac_11_7_io_load),
    .io_mulInput(mac_11_7_io_mulInput),
    .io_addInput(mac_11_7_io_addInput),
    .io_output(mac_11_7_io_output),
    .io_passthrough(mac_11_7_io_passthrough)
  );
  MAC mac_11_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_8_clock),
    .reset(mac_11_8_reset),
    .io_load(mac_11_8_io_load),
    .io_mulInput(mac_11_8_io_mulInput),
    .io_addInput(mac_11_8_io_addInput),
    .io_output(mac_11_8_io_output),
    .io_passthrough(mac_11_8_io_passthrough)
  );
  MAC mac_11_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_9_clock),
    .reset(mac_11_9_reset),
    .io_load(mac_11_9_io_load),
    .io_mulInput(mac_11_9_io_mulInput),
    .io_addInput(mac_11_9_io_addInput),
    .io_output(mac_11_9_io_output),
    .io_passthrough(mac_11_9_io_passthrough)
  );
  MAC mac_11_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_10_clock),
    .reset(mac_11_10_reset),
    .io_load(mac_11_10_io_load),
    .io_mulInput(mac_11_10_io_mulInput),
    .io_addInput(mac_11_10_io_addInput),
    .io_output(mac_11_10_io_output),
    .io_passthrough(mac_11_10_io_passthrough)
  );
  MAC mac_11_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_11_clock),
    .reset(mac_11_11_reset),
    .io_load(mac_11_11_io_load),
    .io_mulInput(mac_11_11_io_mulInput),
    .io_addInput(mac_11_11_io_addInput),
    .io_output(mac_11_11_io_output),
    .io_passthrough(mac_11_11_io_passthrough)
  );
  MAC mac_11_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_12_clock),
    .reset(mac_11_12_reset),
    .io_load(mac_11_12_io_load),
    .io_mulInput(mac_11_12_io_mulInput),
    .io_addInput(mac_11_12_io_addInput),
    .io_output(mac_11_12_io_output),
    .io_passthrough(mac_11_12_io_passthrough)
  );
  MAC mac_11_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_13_clock),
    .reset(mac_11_13_reset),
    .io_load(mac_11_13_io_load),
    .io_mulInput(mac_11_13_io_mulInput),
    .io_addInput(mac_11_13_io_addInput),
    .io_output(mac_11_13_io_output),
    .io_passthrough(mac_11_13_io_passthrough)
  );
  MAC mac_11_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_14_clock),
    .reset(mac_11_14_reset),
    .io_load(mac_11_14_io_load),
    .io_mulInput(mac_11_14_io_mulInput),
    .io_addInput(mac_11_14_io_addInput),
    .io_output(mac_11_14_io_output),
    .io_passthrough(mac_11_14_io_passthrough)
  );
  MAC mac_11_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_15_clock),
    .reset(mac_11_15_reset),
    .io_load(mac_11_15_io_load),
    .io_mulInput(mac_11_15_io_mulInput),
    .io_addInput(mac_11_15_io_addInput),
    .io_output(mac_11_15_io_output),
    .io_passthrough(mac_11_15_io_passthrough)
  );
  MAC mac_11_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_16_clock),
    .reset(mac_11_16_reset),
    .io_load(mac_11_16_io_load),
    .io_mulInput(mac_11_16_io_mulInput),
    .io_addInput(mac_11_16_io_addInput),
    .io_output(mac_11_16_io_output),
    .io_passthrough(mac_11_16_io_passthrough)
  );
  MAC mac_11_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_17_clock),
    .reset(mac_11_17_reset),
    .io_load(mac_11_17_io_load),
    .io_mulInput(mac_11_17_io_mulInput),
    .io_addInput(mac_11_17_io_addInput),
    .io_output(mac_11_17_io_output),
    .io_passthrough(mac_11_17_io_passthrough)
  );
  MAC mac_11_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_18_clock),
    .reset(mac_11_18_reset),
    .io_load(mac_11_18_io_load),
    .io_mulInput(mac_11_18_io_mulInput),
    .io_addInput(mac_11_18_io_addInput),
    .io_output(mac_11_18_io_output),
    .io_passthrough(mac_11_18_io_passthrough)
  );
  MAC mac_11_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_19_clock),
    .reset(mac_11_19_reset),
    .io_load(mac_11_19_io_load),
    .io_mulInput(mac_11_19_io_mulInput),
    .io_addInput(mac_11_19_io_addInput),
    .io_output(mac_11_19_io_output),
    .io_passthrough(mac_11_19_io_passthrough)
  );
  MAC mac_11_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_20_clock),
    .reset(mac_11_20_reset),
    .io_load(mac_11_20_io_load),
    .io_mulInput(mac_11_20_io_mulInput),
    .io_addInput(mac_11_20_io_addInput),
    .io_output(mac_11_20_io_output),
    .io_passthrough(mac_11_20_io_passthrough)
  );
  MAC mac_11_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_21_clock),
    .reset(mac_11_21_reset),
    .io_load(mac_11_21_io_load),
    .io_mulInput(mac_11_21_io_mulInput),
    .io_addInput(mac_11_21_io_addInput),
    .io_output(mac_11_21_io_output),
    .io_passthrough(mac_11_21_io_passthrough)
  );
  MAC mac_11_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_22_clock),
    .reset(mac_11_22_reset),
    .io_load(mac_11_22_io_load),
    .io_mulInput(mac_11_22_io_mulInput),
    .io_addInput(mac_11_22_io_addInput),
    .io_output(mac_11_22_io_output),
    .io_passthrough(mac_11_22_io_passthrough)
  );
  MAC mac_11_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_23_clock),
    .reset(mac_11_23_reset),
    .io_load(mac_11_23_io_load),
    .io_mulInput(mac_11_23_io_mulInput),
    .io_addInput(mac_11_23_io_addInput),
    .io_output(mac_11_23_io_output),
    .io_passthrough(mac_11_23_io_passthrough)
  );
  MAC mac_11_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_24_clock),
    .reset(mac_11_24_reset),
    .io_load(mac_11_24_io_load),
    .io_mulInput(mac_11_24_io_mulInput),
    .io_addInput(mac_11_24_io_addInput),
    .io_output(mac_11_24_io_output),
    .io_passthrough(mac_11_24_io_passthrough)
  );
  MAC mac_11_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_25_clock),
    .reset(mac_11_25_reset),
    .io_load(mac_11_25_io_load),
    .io_mulInput(mac_11_25_io_mulInput),
    .io_addInput(mac_11_25_io_addInput),
    .io_output(mac_11_25_io_output),
    .io_passthrough(mac_11_25_io_passthrough)
  );
  MAC mac_11_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_26_clock),
    .reset(mac_11_26_reset),
    .io_load(mac_11_26_io_load),
    .io_mulInput(mac_11_26_io_mulInput),
    .io_addInput(mac_11_26_io_addInput),
    .io_output(mac_11_26_io_output),
    .io_passthrough(mac_11_26_io_passthrough)
  );
  MAC mac_11_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_27_clock),
    .reset(mac_11_27_reset),
    .io_load(mac_11_27_io_load),
    .io_mulInput(mac_11_27_io_mulInput),
    .io_addInput(mac_11_27_io_addInput),
    .io_output(mac_11_27_io_output),
    .io_passthrough(mac_11_27_io_passthrough)
  );
  MAC mac_11_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_28_clock),
    .reset(mac_11_28_reset),
    .io_load(mac_11_28_io_load),
    .io_mulInput(mac_11_28_io_mulInput),
    .io_addInput(mac_11_28_io_addInput),
    .io_output(mac_11_28_io_output),
    .io_passthrough(mac_11_28_io_passthrough)
  );
  MAC mac_11_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_29_clock),
    .reset(mac_11_29_reset),
    .io_load(mac_11_29_io_load),
    .io_mulInput(mac_11_29_io_mulInput),
    .io_addInput(mac_11_29_io_addInput),
    .io_output(mac_11_29_io_output),
    .io_passthrough(mac_11_29_io_passthrough)
  );
  MAC mac_11_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_30_clock),
    .reset(mac_11_30_reset),
    .io_load(mac_11_30_io_load),
    .io_mulInput(mac_11_30_io_mulInput),
    .io_addInput(mac_11_30_io_addInput),
    .io_output(mac_11_30_io_output),
    .io_passthrough(mac_11_30_io_passthrough)
  );
  MAC mac_11_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_11_31_clock),
    .reset(mac_11_31_reset),
    .io_load(mac_11_31_io_load),
    .io_mulInput(mac_11_31_io_mulInput),
    .io_addInput(mac_11_31_io_addInput),
    .io_output(mac_11_31_io_output),
    .io_passthrough(mac_11_31_io_passthrough)
  );
  MAC mac_12_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_0_clock),
    .reset(mac_12_0_reset),
    .io_load(mac_12_0_io_load),
    .io_mulInput(mac_12_0_io_mulInput),
    .io_addInput(mac_12_0_io_addInput),
    .io_output(mac_12_0_io_output),
    .io_passthrough(mac_12_0_io_passthrough)
  );
  MAC mac_12_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_1_clock),
    .reset(mac_12_1_reset),
    .io_load(mac_12_1_io_load),
    .io_mulInput(mac_12_1_io_mulInput),
    .io_addInput(mac_12_1_io_addInput),
    .io_output(mac_12_1_io_output),
    .io_passthrough(mac_12_1_io_passthrough)
  );
  MAC mac_12_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_2_clock),
    .reset(mac_12_2_reset),
    .io_load(mac_12_2_io_load),
    .io_mulInput(mac_12_2_io_mulInput),
    .io_addInput(mac_12_2_io_addInput),
    .io_output(mac_12_2_io_output),
    .io_passthrough(mac_12_2_io_passthrough)
  );
  MAC mac_12_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_3_clock),
    .reset(mac_12_3_reset),
    .io_load(mac_12_3_io_load),
    .io_mulInput(mac_12_3_io_mulInput),
    .io_addInput(mac_12_3_io_addInput),
    .io_output(mac_12_3_io_output),
    .io_passthrough(mac_12_3_io_passthrough)
  );
  MAC mac_12_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_4_clock),
    .reset(mac_12_4_reset),
    .io_load(mac_12_4_io_load),
    .io_mulInput(mac_12_4_io_mulInput),
    .io_addInput(mac_12_4_io_addInput),
    .io_output(mac_12_4_io_output),
    .io_passthrough(mac_12_4_io_passthrough)
  );
  MAC mac_12_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_5_clock),
    .reset(mac_12_5_reset),
    .io_load(mac_12_5_io_load),
    .io_mulInput(mac_12_5_io_mulInput),
    .io_addInput(mac_12_5_io_addInput),
    .io_output(mac_12_5_io_output),
    .io_passthrough(mac_12_5_io_passthrough)
  );
  MAC mac_12_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_6_clock),
    .reset(mac_12_6_reset),
    .io_load(mac_12_6_io_load),
    .io_mulInput(mac_12_6_io_mulInput),
    .io_addInput(mac_12_6_io_addInput),
    .io_output(mac_12_6_io_output),
    .io_passthrough(mac_12_6_io_passthrough)
  );
  MAC mac_12_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_7_clock),
    .reset(mac_12_7_reset),
    .io_load(mac_12_7_io_load),
    .io_mulInput(mac_12_7_io_mulInput),
    .io_addInput(mac_12_7_io_addInput),
    .io_output(mac_12_7_io_output),
    .io_passthrough(mac_12_7_io_passthrough)
  );
  MAC mac_12_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_8_clock),
    .reset(mac_12_8_reset),
    .io_load(mac_12_8_io_load),
    .io_mulInput(mac_12_8_io_mulInput),
    .io_addInput(mac_12_8_io_addInput),
    .io_output(mac_12_8_io_output),
    .io_passthrough(mac_12_8_io_passthrough)
  );
  MAC mac_12_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_9_clock),
    .reset(mac_12_9_reset),
    .io_load(mac_12_9_io_load),
    .io_mulInput(mac_12_9_io_mulInput),
    .io_addInput(mac_12_9_io_addInput),
    .io_output(mac_12_9_io_output),
    .io_passthrough(mac_12_9_io_passthrough)
  );
  MAC mac_12_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_10_clock),
    .reset(mac_12_10_reset),
    .io_load(mac_12_10_io_load),
    .io_mulInput(mac_12_10_io_mulInput),
    .io_addInput(mac_12_10_io_addInput),
    .io_output(mac_12_10_io_output),
    .io_passthrough(mac_12_10_io_passthrough)
  );
  MAC mac_12_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_11_clock),
    .reset(mac_12_11_reset),
    .io_load(mac_12_11_io_load),
    .io_mulInput(mac_12_11_io_mulInput),
    .io_addInput(mac_12_11_io_addInput),
    .io_output(mac_12_11_io_output),
    .io_passthrough(mac_12_11_io_passthrough)
  );
  MAC mac_12_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_12_clock),
    .reset(mac_12_12_reset),
    .io_load(mac_12_12_io_load),
    .io_mulInput(mac_12_12_io_mulInput),
    .io_addInput(mac_12_12_io_addInput),
    .io_output(mac_12_12_io_output),
    .io_passthrough(mac_12_12_io_passthrough)
  );
  MAC mac_12_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_13_clock),
    .reset(mac_12_13_reset),
    .io_load(mac_12_13_io_load),
    .io_mulInput(mac_12_13_io_mulInput),
    .io_addInput(mac_12_13_io_addInput),
    .io_output(mac_12_13_io_output),
    .io_passthrough(mac_12_13_io_passthrough)
  );
  MAC mac_12_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_14_clock),
    .reset(mac_12_14_reset),
    .io_load(mac_12_14_io_load),
    .io_mulInput(mac_12_14_io_mulInput),
    .io_addInput(mac_12_14_io_addInput),
    .io_output(mac_12_14_io_output),
    .io_passthrough(mac_12_14_io_passthrough)
  );
  MAC mac_12_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_15_clock),
    .reset(mac_12_15_reset),
    .io_load(mac_12_15_io_load),
    .io_mulInput(mac_12_15_io_mulInput),
    .io_addInput(mac_12_15_io_addInput),
    .io_output(mac_12_15_io_output),
    .io_passthrough(mac_12_15_io_passthrough)
  );
  MAC mac_12_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_16_clock),
    .reset(mac_12_16_reset),
    .io_load(mac_12_16_io_load),
    .io_mulInput(mac_12_16_io_mulInput),
    .io_addInput(mac_12_16_io_addInput),
    .io_output(mac_12_16_io_output),
    .io_passthrough(mac_12_16_io_passthrough)
  );
  MAC mac_12_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_17_clock),
    .reset(mac_12_17_reset),
    .io_load(mac_12_17_io_load),
    .io_mulInput(mac_12_17_io_mulInput),
    .io_addInput(mac_12_17_io_addInput),
    .io_output(mac_12_17_io_output),
    .io_passthrough(mac_12_17_io_passthrough)
  );
  MAC mac_12_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_18_clock),
    .reset(mac_12_18_reset),
    .io_load(mac_12_18_io_load),
    .io_mulInput(mac_12_18_io_mulInput),
    .io_addInput(mac_12_18_io_addInput),
    .io_output(mac_12_18_io_output),
    .io_passthrough(mac_12_18_io_passthrough)
  );
  MAC mac_12_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_19_clock),
    .reset(mac_12_19_reset),
    .io_load(mac_12_19_io_load),
    .io_mulInput(mac_12_19_io_mulInput),
    .io_addInput(mac_12_19_io_addInput),
    .io_output(mac_12_19_io_output),
    .io_passthrough(mac_12_19_io_passthrough)
  );
  MAC mac_12_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_20_clock),
    .reset(mac_12_20_reset),
    .io_load(mac_12_20_io_load),
    .io_mulInput(mac_12_20_io_mulInput),
    .io_addInput(mac_12_20_io_addInput),
    .io_output(mac_12_20_io_output),
    .io_passthrough(mac_12_20_io_passthrough)
  );
  MAC mac_12_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_21_clock),
    .reset(mac_12_21_reset),
    .io_load(mac_12_21_io_load),
    .io_mulInput(mac_12_21_io_mulInput),
    .io_addInput(mac_12_21_io_addInput),
    .io_output(mac_12_21_io_output),
    .io_passthrough(mac_12_21_io_passthrough)
  );
  MAC mac_12_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_22_clock),
    .reset(mac_12_22_reset),
    .io_load(mac_12_22_io_load),
    .io_mulInput(mac_12_22_io_mulInput),
    .io_addInput(mac_12_22_io_addInput),
    .io_output(mac_12_22_io_output),
    .io_passthrough(mac_12_22_io_passthrough)
  );
  MAC mac_12_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_23_clock),
    .reset(mac_12_23_reset),
    .io_load(mac_12_23_io_load),
    .io_mulInput(mac_12_23_io_mulInput),
    .io_addInput(mac_12_23_io_addInput),
    .io_output(mac_12_23_io_output),
    .io_passthrough(mac_12_23_io_passthrough)
  );
  MAC mac_12_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_24_clock),
    .reset(mac_12_24_reset),
    .io_load(mac_12_24_io_load),
    .io_mulInput(mac_12_24_io_mulInput),
    .io_addInput(mac_12_24_io_addInput),
    .io_output(mac_12_24_io_output),
    .io_passthrough(mac_12_24_io_passthrough)
  );
  MAC mac_12_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_25_clock),
    .reset(mac_12_25_reset),
    .io_load(mac_12_25_io_load),
    .io_mulInput(mac_12_25_io_mulInput),
    .io_addInput(mac_12_25_io_addInput),
    .io_output(mac_12_25_io_output),
    .io_passthrough(mac_12_25_io_passthrough)
  );
  MAC mac_12_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_26_clock),
    .reset(mac_12_26_reset),
    .io_load(mac_12_26_io_load),
    .io_mulInput(mac_12_26_io_mulInput),
    .io_addInput(mac_12_26_io_addInput),
    .io_output(mac_12_26_io_output),
    .io_passthrough(mac_12_26_io_passthrough)
  );
  MAC mac_12_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_27_clock),
    .reset(mac_12_27_reset),
    .io_load(mac_12_27_io_load),
    .io_mulInput(mac_12_27_io_mulInput),
    .io_addInput(mac_12_27_io_addInput),
    .io_output(mac_12_27_io_output),
    .io_passthrough(mac_12_27_io_passthrough)
  );
  MAC mac_12_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_28_clock),
    .reset(mac_12_28_reset),
    .io_load(mac_12_28_io_load),
    .io_mulInput(mac_12_28_io_mulInput),
    .io_addInput(mac_12_28_io_addInput),
    .io_output(mac_12_28_io_output),
    .io_passthrough(mac_12_28_io_passthrough)
  );
  MAC mac_12_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_29_clock),
    .reset(mac_12_29_reset),
    .io_load(mac_12_29_io_load),
    .io_mulInput(mac_12_29_io_mulInput),
    .io_addInput(mac_12_29_io_addInput),
    .io_output(mac_12_29_io_output),
    .io_passthrough(mac_12_29_io_passthrough)
  );
  MAC mac_12_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_30_clock),
    .reset(mac_12_30_reset),
    .io_load(mac_12_30_io_load),
    .io_mulInput(mac_12_30_io_mulInput),
    .io_addInput(mac_12_30_io_addInput),
    .io_output(mac_12_30_io_output),
    .io_passthrough(mac_12_30_io_passthrough)
  );
  MAC mac_12_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_12_31_clock),
    .reset(mac_12_31_reset),
    .io_load(mac_12_31_io_load),
    .io_mulInput(mac_12_31_io_mulInput),
    .io_addInput(mac_12_31_io_addInput),
    .io_output(mac_12_31_io_output),
    .io_passthrough(mac_12_31_io_passthrough)
  );
  MAC mac_13_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_0_clock),
    .reset(mac_13_0_reset),
    .io_load(mac_13_0_io_load),
    .io_mulInput(mac_13_0_io_mulInput),
    .io_addInput(mac_13_0_io_addInput),
    .io_output(mac_13_0_io_output),
    .io_passthrough(mac_13_0_io_passthrough)
  );
  MAC mac_13_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_1_clock),
    .reset(mac_13_1_reset),
    .io_load(mac_13_1_io_load),
    .io_mulInput(mac_13_1_io_mulInput),
    .io_addInput(mac_13_1_io_addInput),
    .io_output(mac_13_1_io_output),
    .io_passthrough(mac_13_1_io_passthrough)
  );
  MAC mac_13_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_2_clock),
    .reset(mac_13_2_reset),
    .io_load(mac_13_2_io_load),
    .io_mulInput(mac_13_2_io_mulInput),
    .io_addInput(mac_13_2_io_addInput),
    .io_output(mac_13_2_io_output),
    .io_passthrough(mac_13_2_io_passthrough)
  );
  MAC mac_13_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_3_clock),
    .reset(mac_13_3_reset),
    .io_load(mac_13_3_io_load),
    .io_mulInput(mac_13_3_io_mulInput),
    .io_addInput(mac_13_3_io_addInput),
    .io_output(mac_13_3_io_output),
    .io_passthrough(mac_13_3_io_passthrough)
  );
  MAC mac_13_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_4_clock),
    .reset(mac_13_4_reset),
    .io_load(mac_13_4_io_load),
    .io_mulInput(mac_13_4_io_mulInput),
    .io_addInput(mac_13_4_io_addInput),
    .io_output(mac_13_4_io_output),
    .io_passthrough(mac_13_4_io_passthrough)
  );
  MAC mac_13_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_5_clock),
    .reset(mac_13_5_reset),
    .io_load(mac_13_5_io_load),
    .io_mulInput(mac_13_5_io_mulInput),
    .io_addInput(mac_13_5_io_addInput),
    .io_output(mac_13_5_io_output),
    .io_passthrough(mac_13_5_io_passthrough)
  );
  MAC mac_13_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_6_clock),
    .reset(mac_13_6_reset),
    .io_load(mac_13_6_io_load),
    .io_mulInput(mac_13_6_io_mulInput),
    .io_addInput(mac_13_6_io_addInput),
    .io_output(mac_13_6_io_output),
    .io_passthrough(mac_13_6_io_passthrough)
  );
  MAC mac_13_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_7_clock),
    .reset(mac_13_7_reset),
    .io_load(mac_13_7_io_load),
    .io_mulInput(mac_13_7_io_mulInput),
    .io_addInput(mac_13_7_io_addInput),
    .io_output(mac_13_7_io_output),
    .io_passthrough(mac_13_7_io_passthrough)
  );
  MAC mac_13_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_8_clock),
    .reset(mac_13_8_reset),
    .io_load(mac_13_8_io_load),
    .io_mulInput(mac_13_8_io_mulInput),
    .io_addInput(mac_13_8_io_addInput),
    .io_output(mac_13_8_io_output),
    .io_passthrough(mac_13_8_io_passthrough)
  );
  MAC mac_13_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_9_clock),
    .reset(mac_13_9_reset),
    .io_load(mac_13_9_io_load),
    .io_mulInput(mac_13_9_io_mulInput),
    .io_addInput(mac_13_9_io_addInput),
    .io_output(mac_13_9_io_output),
    .io_passthrough(mac_13_9_io_passthrough)
  );
  MAC mac_13_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_10_clock),
    .reset(mac_13_10_reset),
    .io_load(mac_13_10_io_load),
    .io_mulInput(mac_13_10_io_mulInput),
    .io_addInput(mac_13_10_io_addInput),
    .io_output(mac_13_10_io_output),
    .io_passthrough(mac_13_10_io_passthrough)
  );
  MAC mac_13_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_11_clock),
    .reset(mac_13_11_reset),
    .io_load(mac_13_11_io_load),
    .io_mulInput(mac_13_11_io_mulInput),
    .io_addInput(mac_13_11_io_addInput),
    .io_output(mac_13_11_io_output),
    .io_passthrough(mac_13_11_io_passthrough)
  );
  MAC mac_13_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_12_clock),
    .reset(mac_13_12_reset),
    .io_load(mac_13_12_io_load),
    .io_mulInput(mac_13_12_io_mulInput),
    .io_addInput(mac_13_12_io_addInput),
    .io_output(mac_13_12_io_output),
    .io_passthrough(mac_13_12_io_passthrough)
  );
  MAC mac_13_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_13_clock),
    .reset(mac_13_13_reset),
    .io_load(mac_13_13_io_load),
    .io_mulInput(mac_13_13_io_mulInput),
    .io_addInput(mac_13_13_io_addInput),
    .io_output(mac_13_13_io_output),
    .io_passthrough(mac_13_13_io_passthrough)
  );
  MAC mac_13_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_14_clock),
    .reset(mac_13_14_reset),
    .io_load(mac_13_14_io_load),
    .io_mulInput(mac_13_14_io_mulInput),
    .io_addInput(mac_13_14_io_addInput),
    .io_output(mac_13_14_io_output),
    .io_passthrough(mac_13_14_io_passthrough)
  );
  MAC mac_13_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_15_clock),
    .reset(mac_13_15_reset),
    .io_load(mac_13_15_io_load),
    .io_mulInput(mac_13_15_io_mulInput),
    .io_addInput(mac_13_15_io_addInput),
    .io_output(mac_13_15_io_output),
    .io_passthrough(mac_13_15_io_passthrough)
  );
  MAC mac_13_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_16_clock),
    .reset(mac_13_16_reset),
    .io_load(mac_13_16_io_load),
    .io_mulInput(mac_13_16_io_mulInput),
    .io_addInput(mac_13_16_io_addInput),
    .io_output(mac_13_16_io_output),
    .io_passthrough(mac_13_16_io_passthrough)
  );
  MAC mac_13_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_17_clock),
    .reset(mac_13_17_reset),
    .io_load(mac_13_17_io_load),
    .io_mulInput(mac_13_17_io_mulInput),
    .io_addInput(mac_13_17_io_addInput),
    .io_output(mac_13_17_io_output),
    .io_passthrough(mac_13_17_io_passthrough)
  );
  MAC mac_13_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_18_clock),
    .reset(mac_13_18_reset),
    .io_load(mac_13_18_io_load),
    .io_mulInput(mac_13_18_io_mulInput),
    .io_addInput(mac_13_18_io_addInput),
    .io_output(mac_13_18_io_output),
    .io_passthrough(mac_13_18_io_passthrough)
  );
  MAC mac_13_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_19_clock),
    .reset(mac_13_19_reset),
    .io_load(mac_13_19_io_load),
    .io_mulInput(mac_13_19_io_mulInput),
    .io_addInput(mac_13_19_io_addInput),
    .io_output(mac_13_19_io_output),
    .io_passthrough(mac_13_19_io_passthrough)
  );
  MAC mac_13_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_20_clock),
    .reset(mac_13_20_reset),
    .io_load(mac_13_20_io_load),
    .io_mulInput(mac_13_20_io_mulInput),
    .io_addInput(mac_13_20_io_addInput),
    .io_output(mac_13_20_io_output),
    .io_passthrough(mac_13_20_io_passthrough)
  );
  MAC mac_13_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_21_clock),
    .reset(mac_13_21_reset),
    .io_load(mac_13_21_io_load),
    .io_mulInput(mac_13_21_io_mulInput),
    .io_addInput(mac_13_21_io_addInput),
    .io_output(mac_13_21_io_output),
    .io_passthrough(mac_13_21_io_passthrough)
  );
  MAC mac_13_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_22_clock),
    .reset(mac_13_22_reset),
    .io_load(mac_13_22_io_load),
    .io_mulInput(mac_13_22_io_mulInput),
    .io_addInput(mac_13_22_io_addInput),
    .io_output(mac_13_22_io_output),
    .io_passthrough(mac_13_22_io_passthrough)
  );
  MAC mac_13_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_23_clock),
    .reset(mac_13_23_reset),
    .io_load(mac_13_23_io_load),
    .io_mulInput(mac_13_23_io_mulInput),
    .io_addInput(mac_13_23_io_addInput),
    .io_output(mac_13_23_io_output),
    .io_passthrough(mac_13_23_io_passthrough)
  );
  MAC mac_13_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_24_clock),
    .reset(mac_13_24_reset),
    .io_load(mac_13_24_io_load),
    .io_mulInput(mac_13_24_io_mulInput),
    .io_addInput(mac_13_24_io_addInput),
    .io_output(mac_13_24_io_output),
    .io_passthrough(mac_13_24_io_passthrough)
  );
  MAC mac_13_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_25_clock),
    .reset(mac_13_25_reset),
    .io_load(mac_13_25_io_load),
    .io_mulInput(mac_13_25_io_mulInput),
    .io_addInput(mac_13_25_io_addInput),
    .io_output(mac_13_25_io_output),
    .io_passthrough(mac_13_25_io_passthrough)
  );
  MAC mac_13_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_26_clock),
    .reset(mac_13_26_reset),
    .io_load(mac_13_26_io_load),
    .io_mulInput(mac_13_26_io_mulInput),
    .io_addInput(mac_13_26_io_addInput),
    .io_output(mac_13_26_io_output),
    .io_passthrough(mac_13_26_io_passthrough)
  );
  MAC mac_13_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_27_clock),
    .reset(mac_13_27_reset),
    .io_load(mac_13_27_io_load),
    .io_mulInput(mac_13_27_io_mulInput),
    .io_addInput(mac_13_27_io_addInput),
    .io_output(mac_13_27_io_output),
    .io_passthrough(mac_13_27_io_passthrough)
  );
  MAC mac_13_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_28_clock),
    .reset(mac_13_28_reset),
    .io_load(mac_13_28_io_load),
    .io_mulInput(mac_13_28_io_mulInput),
    .io_addInput(mac_13_28_io_addInput),
    .io_output(mac_13_28_io_output),
    .io_passthrough(mac_13_28_io_passthrough)
  );
  MAC mac_13_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_29_clock),
    .reset(mac_13_29_reset),
    .io_load(mac_13_29_io_load),
    .io_mulInput(mac_13_29_io_mulInput),
    .io_addInput(mac_13_29_io_addInput),
    .io_output(mac_13_29_io_output),
    .io_passthrough(mac_13_29_io_passthrough)
  );
  MAC mac_13_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_30_clock),
    .reset(mac_13_30_reset),
    .io_load(mac_13_30_io_load),
    .io_mulInput(mac_13_30_io_mulInput),
    .io_addInput(mac_13_30_io_addInput),
    .io_output(mac_13_30_io_output),
    .io_passthrough(mac_13_30_io_passthrough)
  );
  MAC mac_13_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_13_31_clock),
    .reset(mac_13_31_reset),
    .io_load(mac_13_31_io_load),
    .io_mulInput(mac_13_31_io_mulInput),
    .io_addInput(mac_13_31_io_addInput),
    .io_output(mac_13_31_io_output),
    .io_passthrough(mac_13_31_io_passthrough)
  );
  MAC mac_14_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_0_clock),
    .reset(mac_14_0_reset),
    .io_load(mac_14_0_io_load),
    .io_mulInput(mac_14_0_io_mulInput),
    .io_addInput(mac_14_0_io_addInput),
    .io_output(mac_14_0_io_output),
    .io_passthrough(mac_14_0_io_passthrough)
  );
  MAC mac_14_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_1_clock),
    .reset(mac_14_1_reset),
    .io_load(mac_14_1_io_load),
    .io_mulInput(mac_14_1_io_mulInput),
    .io_addInput(mac_14_1_io_addInput),
    .io_output(mac_14_1_io_output),
    .io_passthrough(mac_14_1_io_passthrough)
  );
  MAC mac_14_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_2_clock),
    .reset(mac_14_2_reset),
    .io_load(mac_14_2_io_load),
    .io_mulInput(mac_14_2_io_mulInput),
    .io_addInput(mac_14_2_io_addInput),
    .io_output(mac_14_2_io_output),
    .io_passthrough(mac_14_2_io_passthrough)
  );
  MAC mac_14_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_3_clock),
    .reset(mac_14_3_reset),
    .io_load(mac_14_3_io_load),
    .io_mulInput(mac_14_3_io_mulInput),
    .io_addInput(mac_14_3_io_addInput),
    .io_output(mac_14_3_io_output),
    .io_passthrough(mac_14_3_io_passthrough)
  );
  MAC mac_14_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_4_clock),
    .reset(mac_14_4_reset),
    .io_load(mac_14_4_io_load),
    .io_mulInput(mac_14_4_io_mulInput),
    .io_addInput(mac_14_4_io_addInput),
    .io_output(mac_14_4_io_output),
    .io_passthrough(mac_14_4_io_passthrough)
  );
  MAC mac_14_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_5_clock),
    .reset(mac_14_5_reset),
    .io_load(mac_14_5_io_load),
    .io_mulInput(mac_14_5_io_mulInput),
    .io_addInput(mac_14_5_io_addInput),
    .io_output(mac_14_5_io_output),
    .io_passthrough(mac_14_5_io_passthrough)
  );
  MAC mac_14_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_6_clock),
    .reset(mac_14_6_reset),
    .io_load(mac_14_6_io_load),
    .io_mulInput(mac_14_6_io_mulInput),
    .io_addInput(mac_14_6_io_addInput),
    .io_output(mac_14_6_io_output),
    .io_passthrough(mac_14_6_io_passthrough)
  );
  MAC mac_14_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_7_clock),
    .reset(mac_14_7_reset),
    .io_load(mac_14_7_io_load),
    .io_mulInput(mac_14_7_io_mulInput),
    .io_addInput(mac_14_7_io_addInput),
    .io_output(mac_14_7_io_output),
    .io_passthrough(mac_14_7_io_passthrough)
  );
  MAC mac_14_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_8_clock),
    .reset(mac_14_8_reset),
    .io_load(mac_14_8_io_load),
    .io_mulInput(mac_14_8_io_mulInput),
    .io_addInput(mac_14_8_io_addInput),
    .io_output(mac_14_8_io_output),
    .io_passthrough(mac_14_8_io_passthrough)
  );
  MAC mac_14_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_9_clock),
    .reset(mac_14_9_reset),
    .io_load(mac_14_9_io_load),
    .io_mulInput(mac_14_9_io_mulInput),
    .io_addInput(mac_14_9_io_addInput),
    .io_output(mac_14_9_io_output),
    .io_passthrough(mac_14_9_io_passthrough)
  );
  MAC mac_14_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_10_clock),
    .reset(mac_14_10_reset),
    .io_load(mac_14_10_io_load),
    .io_mulInput(mac_14_10_io_mulInput),
    .io_addInput(mac_14_10_io_addInput),
    .io_output(mac_14_10_io_output),
    .io_passthrough(mac_14_10_io_passthrough)
  );
  MAC mac_14_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_11_clock),
    .reset(mac_14_11_reset),
    .io_load(mac_14_11_io_load),
    .io_mulInput(mac_14_11_io_mulInput),
    .io_addInput(mac_14_11_io_addInput),
    .io_output(mac_14_11_io_output),
    .io_passthrough(mac_14_11_io_passthrough)
  );
  MAC mac_14_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_12_clock),
    .reset(mac_14_12_reset),
    .io_load(mac_14_12_io_load),
    .io_mulInput(mac_14_12_io_mulInput),
    .io_addInput(mac_14_12_io_addInput),
    .io_output(mac_14_12_io_output),
    .io_passthrough(mac_14_12_io_passthrough)
  );
  MAC mac_14_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_13_clock),
    .reset(mac_14_13_reset),
    .io_load(mac_14_13_io_load),
    .io_mulInput(mac_14_13_io_mulInput),
    .io_addInput(mac_14_13_io_addInput),
    .io_output(mac_14_13_io_output),
    .io_passthrough(mac_14_13_io_passthrough)
  );
  MAC mac_14_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_14_clock),
    .reset(mac_14_14_reset),
    .io_load(mac_14_14_io_load),
    .io_mulInput(mac_14_14_io_mulInput),
    .io_addInput(mac_14_14_io_addInput),
    .io_output(mac_14_14_io_output),
    .io_passthrough(mac_14_14_io_passthrough)
  );
  MAC mac_14_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_15_clock),
    .reset(mac_14_15_reset),
    .io_load(mac_14_15_io_load),
    .io_mulInput(mac_14_15_io_mulInput),
    .io_addInput(mac_14_15_io_addInput),
    .io_output(mac_14_15_io_output),
    .io_passthrough(mac_14_15_io_passthrough)
  );
  MAC mac_14_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_16_clock),
    .reset(mac_14_16_reset),
    .io_load(mac_14_16_io_load),
    .io_mulInput(mac_14_16_io_mulInput),
    .io_addInput(mac_14_16_io_addInput),
    .io_output(mac_14_16_io_output),
    .io_passthrough(mac_14_16_io_passthrough)
  );
  MAC mac_14_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_17_clock),
    .reset(mac_14_17_reset),
    .io_load(mac_14_17_io_load),
    .io_mulInput(mac_14_17_io_mulInput),
    .io_addInput(mac_14_17_io_addInput),
    .io_output(mac_14_17_io_output),
    .io_passthrough(mac_14_17_io_passthrough)
  );
  MAC mac_14_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_18_clock),
    .reset(mac_14_18_reset),
    .io_load(mac_14_18_io_load),
    .io_mulInput(mac_14_18_io_mulInput),
    .io_addInput(mac_14_18_io_addInput),
    .io_output(mac_14_18_io_output),
    .io_passthrough(mac_14_18_io_passthrough)
  );
  MAC mac_14_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_19_clock),
    .reset(mac_14_19_reset),
    .io_load(mac_14_19_io_load),
    .io_mulInput(mac_14_19_io_mulInput),
    .io_addInput(mac_14_19_io_addInput),
    .io_output(mac_14_19_io_output),
    .io_passthrough(mac_14_19_io_passthrough)
  );
  MAC mac_14_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_20_clock),
    .reset(mac_14_20_reset),
    .io_load(mac_14_20_io_load),
    .io_mulInput(mac_14_20_io_mulInput),
    .io_addInput(mac_14_20_io_addInput),
    .io_output(mac_14_20_io_output),
    .io_passthrough(mac_14_20_io_passthrough)
  );
  MAC mac_14_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_21_clock),
    .reset(mac_14_21_reset),
    .io_load(mac_14_21_io_load),
    .io_mulInput(mac_14_21_io_mulInput),
    .io_addInput(mac_14_21_io_addInput),
    .io_output(mac_14_21_io_output),
    .io_passthrough(mac_14_21_io_passthrough)
  );
  MAC mac_14_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_22_clock),
    .reset(mac_14_22_reset),
    .io_load(mac_14_22_io_load),
    .io_mulInput(mac_14_22_io_mulInput),
    .io_addInput(mac_14_22_io_addInput),
    .io_output(mac_14_22_io_output),
    .io_passthrough(mac_14_22_io_passthrough)
  );
  MAC mac_14_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_23_clock),
    .reset(mac_14_23_reset),
    .io_load(mac_14_23_io_load),
    .io_mulInput(mac_14_23_io_mulInput),
    .io_addInput(mac_14_23_io_addInput),
    .io_output(mac_14_23_io_output),
    .io_passthrough(mac_14_23_io_passthrough)
  );
  MAC mac_14_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_24_clock),
    .reset(mac_14_24_reset),
    .io_load(mac_14_24_io_load),
    .io_mulInput(mac_14_24_io_mulInput),
    .io_addInput(mac_14_24_io_addInput),
    .io_output(mac_14_24_io_output),
    .io_passthrough(mac_14_24_io_passthrough)
  );
  MAC mac_14_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_25_clock),
    .reset(mac_14_25_reset),
    .io_load(mac_14_25_io_load),
    .io_mulInput(mac_14_25_io_mulInput),
    .io_addInput(mac_14_25_io_addInput),
    .io_output(mac_14_25_io_output),
    .io_passthrough(mac_14_25_io_passthrough)
  );
  MAC mac_14_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_26_clock),
    .reset(mac_14_26_reset),
    .io_load(mac_14_26_io_load),
    .io_mulInput(mac_14_26_io_mulInput),
    .io_addInput(mac_14_26_io_addInput),
    .io_output(mac_14_26_io_output),
    .io_passthrough(mac_14_26_io_passthrough)
  );
  MAC mac_14_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_27_clock),
    .reset(mac_14_27_reset),
    .io_load(mac_14_27_io_load),
    .io_mulInput(mac_14_27_io_mulInput),
    .io_addInput(mac_14_27_io_addInput),
    .io_output(mac_14_27_io_output),
    .io_passthrough(mac_14_27_io_passthrough)
  );
  MAC mac_14_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_28_clock),
    .reset(mac_14_28_reset),
    .io_load(mac_14_28_io_load),
    .io_mulInput(mac_14_28_io_mulInput),
    .io_addInput(mac_14_28_io_addInput),
    .io_output(mac_14_28_io_output),
    .io_passthrough(mac_14_28_io_passthrough)
  );
  MAC mac_14_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_29_clock),
    .reset(mac_14_29_reset),
    .io_load(mac_14_29_io_load),
    .io_mulInput(mac_14_29_io_mulInput),
    .io_addInput(mac_14_29_io_addInput),
    .io_output(mac_14_29_io_output),
    .io_passthrough(mac_14_29_io_passthrough)
  );
  MAC mac_14_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_30_clock),
    .reset(mac_14_30_reset),
    .io_load(mac_14_30_io_load),
    .io_mulInput(mac_14_30_io_mulInput),
    .io_addInput(mac_14_30_io_addInput),
    .io_output(mac_14_30_io_output),
    .io_passthrough(mac_14_30_io_passthrough)
  );
  MAC mac_14_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_14_31_clock),
    .reset(mac_14_31_reset),
    .io_load(mac_14_31_io_load),
    .io_mulInput(mac_14_31_io_mulInput),
    .io_addInput(mac_14_31_io_addInput),
    .io_output(mac_14_31_io_output),
    .io_passthrough(mac_14_31_io_passthrough)
  );
  MAC mac_15_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_0_clock),
    .reset(mac_15_0_reset),
    .io_load(mac_15_0_io_load),
    .io_mulInput(mac_15_0_io_mulInput),
    .io_addInput(mac_15_0_io_addInput),
    .io_output(mac_15_0_io_output),
    .io_passthrough(mac_15_0_io_passthrough)
  );
  MAC mac_15_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_1_clock),
    .reset(mac_15_1_reset),
    .io_load(mac_15_1_io_load),
    .io_mulInput(mac_15_1_io_mulInput),
    .io_addInput(mac_15_1_io_addInput),
    .io_output(mac_15_1_io_output),
    .io_passthrough(mac_15_1_io_passthrough)
  );
  MAC mac_15_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_2_clock),
    .reset(mac_15_2_reset),
    .io_load(mac_15_2_io_load),
    .io_mulInput(mac_15_2_io_mulInput),
    .io_addInput(mac_15_2_io_addInput),
    .io_output(mac_15_2_io_output),
    .io_passthrough(mac_15_2_io_passthrough)
  );
  MAC mac_15_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_3_clock),
    .reset(mac_15_3_reset),
    .io_load(mac_15_3_io_load),
    .io_mulInput(mac_15_3_io_mulInput),
    .io_addInput(mac_15_3_io_addInput),
    .io_output(mac_15_3_io_output),
    .io_passthrough(mac_15_3_io_passthrough)
  );
  MAC mac_15_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_4_clock),
    .reset(mac_15_4_reset),
    .io_load(mac_15_4_io_load),
    .io_mulInput(mac_15_4_io_mulInput),
    .io_addInput(mac_15_4_io_addInput),
    .io_output(mac_15_4_io_output),
    .io_passthrough(mac_15_4_io_passthrough)
  );
  MAC mac_15_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_5_clock),
    .reset(mac_15_5_reset),
    .io_load(mac_15_5_io_load),
    .io_mulInput(mac_15_5_io_mulInput),
    .io_addInput(mac_15_5_io_addInput),
    .io_output(mac_15_5_io_output),
    .io_passthrough(mac_15_5_io_passthrough)
  );
  MAC mac_15_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_6_clock),
    .reset(mac_15_6_reset),
    .io_load(mac_15_6_io_load),
    .io_mulInput(mac_15_6_io_mulInput),
    .io_addInput(mac_15_6_io_addInput),
    .io_output(mac_15_6_io_output),
    .io_passthrough(mac_15_6_io_passthrough)
  );
  MAC mac_15_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_7_clock),
    .reset(mac_15_7_reset),
    .io_load(mac_15_7_io_load),
    .io_mulInput(mac_15_7_io_mulInput),
    .io_addInput(mac_15_7_io_addInput),
    .io_output(mac_15_7_io_output),
    .io_passthrough(mac_15_7_io_passthrough)
  );
  MAC mac_15_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_8_clock),
    .reset(mac_15_8_reset),
    .io_load(mac_15_8_io_load),
    .io_mulInput(mac_15_8_io_mulInput),
    .io_addInput(mac_15_8_io_addInput),
    .io_output(mac_15_8_io_output),
    .io_passthrough(mac_15_8_io_passthrough)
  );
  MAC mac_15_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_9_clock),
    .reset(mac_15_9_reset),
    .io_load(mac_15_9_io_load),
    .io_mulInput(mac_15_9_io_mulInput),
    .io_addInput(mac_15_9_io_addInput),
    .io_output(mac_15_9_io_output),
    .io_passthrough(mac_15_9_io_passthrough)
  );
  MAC mac_15_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_10_clock),
    .reset(mac_15_10_reset),
    .io_load(mac_15_10_io_load),
    .io_mulInput(mac_15_10_io_mulInput),
    .io_addInput(mac_15_10_io_addInput),
    .io_output(mac_15_10_io_output),
    .io_passthrough(mac_15_10_io_passthrough)
  );
  MAC mac_15_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_11_clock),
    .reset(mac_15_11_reset),
    .io_load(mac_15_11_io_load),
    .io_mulInput(mac_15_11_io_mulInput),
    .io_addInput(mac_15_11_io_addInput),
    .io_output(mac_15_11_io_output),
    .io_passthrough(mac_15_11_io_passthrough)
  );
  MAC mac_15_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_12_clock),
    .reset(mac_15_12_reset),
    .io_load(mac_15_12_io_load),
    .io_mulInput(mac_15_12_io_mulInput),
    .io_addInput(mac_15_12_io_addInput),
    .io_output(mac_15_12_io_output),
    .io_passthrough(mac_15_12_io_passthrough)
  );
  MAC mac_15_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_13_clock),
    .reset(mac_15_13_reset),
    .io_load(mac_15_13_io_load),
    .io_mulInput(mac_15_13_io_mulInput),
    .io_addInput(mac_15_13_io_addInput),
    .io_output(mac_15_13_io_output),
    .io_passthrough(mac_15_13_io_passthrough)
  );
  MAC mac_15_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_14_clock),
    .reset(mac_15_14_reset),
    .io_load(mac_15_14_io_load),
    .io_mulInput(mac_15_14_io_mulInput),
    .io_addInput(mac_15_14_io_addInput),
    .io_output(mac_15_14_io_output),
    .io_passthrough(mac_15_14_io_passthrough)
  );
  MAC mac_15_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_15_clock),
    .reset(mac_15_15_reset),
    .io_load(mac_15_15_io_load),
    .io_mulInput(mac_15_15_io_mulInput),
    .io_addInput(mac_15_15_io_addInput),
    .io_output(mac_15_15_io_output),
    .io_passthrough(mac_15_15_io_passthrough)
  );
  MAC mac_15_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_16_clock),
    .reset(mac_15_16_reset),
    .io_load(mac_15_16_io_load),
    .io_mulInput(mac_15_16_io_mulInput),
    .io_addInput(mac_15_16_io_addInput),
    .io_output(mac_15_16_io_output),
    .io_passthrough(mac_15_16_io_passthrough)
  );
  MAC mac_15_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_17_clock),
    .reset(mac_15_17_reset),
    .io_load(mac_15_17_io_load),
    .io_mulInput(mac_15_17_io_mulInput),
    .io_addInput(mac_15_17_io_addInput),
    .io_output(mac_15_17_io_output),
    .io_passthrough(mac_15_17_io_passthrough)
  );
  MAC mac_15_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_18_clock),
    .reset(mac_15_18_reset),
    .io_load(mac_15_18_io_load),
    .io_mulInput(mac_15_18_io_mulInput),
    .io_addInput(mac_15_18_io_addInput),
    .io_output(mac_15_18_io_output),
    .io_passthrough(mac_15_18_io_passthrough)
  );
  MAC mac_15_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_19_clock),
    .reset(mac_15_19_reset),
    .io_load(mac_15_19_io_load),
    .io_mulInput(mac_15_19_io_mulInput),
    .io_addInput(mac_15_19_io_addInput),
    .io_output(mac_15_19_io_output),
    .io_passthrough(mac_15_19_io_passthrough)
  );
  MAC mac_15_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_20_clock),
    .reset(mac_15_20_reset),
    .io_load(mac_15_20_io_load),
    .io_mulInput(mac_15_20_io_mulInput),
    .io_addInput(mac_15_20_io_addInput),
    .io_output(mac_15_20_io_output),
    .io_passthrough(mac_15_20_io_passthrough)
  );
  MAC mac_15_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_21_clock),
    .reset(mac_15_21_reset),
    .io_load(mac_15_21_io_load),
    .io_mulInput(mac_15_21_io_mulInput),
    .io_addInput(mac_15_21_io_addInput),
    .io_output(mac_15_21_io_output),
    .io_passthrough(mac_15_21_io_passthrough)
  );
  MAC mac_15_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_22_clock),
    .reset(mac_15_22_reset),
    .io_load(mac_15_22_io_load),
    .io_mulInput(mac_15_22_io_mulInput),
    .io_addInput(mac_15_22_io_addInput),
    .io_output(mac_15_22_io_output),
    .io_passthrough(mac_15_22_io_passthrough)
  );
  MAC mac_15_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_23_clock),
    .reset(mac_15_23_reset),
    .io_load(mac_15_23_io_load),
    .io_mulInput(mac_15_23_io_mulInput),
    .io_addInput(mac_15_23_io_addInput),
    .io_output(mac_15_23_io_output),
    .io_passthrough(mac_15_23_io_passthrough)
  );
  MAC mac_15_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_24_clock),
    .reset(mac_15_24_reset),
    .io_load(mac_15_24_io_load),
    .io_mulInput(mac_15_24_io_mulInput),
    .io_addInput(mac_15_24_io_addInput),
    .io_output(mac_15_24_io_output),
    .io_passthrough(mac_15_24_io_passthrough)
  );
  MAC mac_15_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_25_clock),
    .reset(mac_15_25_reset),
    .io_load(mac_15_25_io_load),
    .io_mulInput(mac_15_25_io_mulInput),
    .io_addInput(mac_15_25_io_addInput),
    .io_output(mac_15_25_io_output),
    .io_passthrough(mac_15_25_io_passthrough)
  );
  MAC mac_15_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_26_clock),
    .reset(mac_15_26_reset),
    .io_load(mac_15_26_io_load),
    .io_mulInput(mac_15_26_io_mulInput),
    .io_addInput(mac_15_26_io_addInput),
    .io_output(mac_15_26_io_output),
    .io_passthrough(mac_15_26_io_passthrough)
  );
  MAC mac_15_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_27_clock),
    .reset(mac_15_27_reset),
    .io_load(mac_15_27_io_load),
    .io_mulInput(mac_15_27_io_mulInput),
    .io_addInput(mac_15_27_io_addInput),
    .io_output(mac_15_27_io_output),
    .io_passthrough(mac_15_27_io_passthrough)
  );
  MAC mac_15_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_28_clock),
    .reset(mac_15_28_reset),
    .io_load(mac_15_28_io_load),
    .io_mulInput(mac_15_28_io_mulInput),
    .io_addInput(mac_15_28_io_addInput),
    .io_output(mac_15_28_io_output),
    .io_passthrough(mac_15_28_io_passthrough)
  );
  MAC mac_15_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_29_clock),
    .reset(mac_15_29_reset),
    .io_load(mac_15_29_io_load),
    .io_mulInput(mac_15_29_io_mulInput),
    .io_addInput(mac_15_29_io_addInput),
    .io_output(mac_15_29_io_output),
    .io_passthrough(mac_15_29_io_passthrough)
  );
  MAC mac_15_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_30_clock),
    .reset(mac_15_30_reset),
    .io_load(mac_15_30_io_load),
    .io_mulInput(mac_15_30_io_mulInput),
    .io_addInput(mac_15_30_io_addInput),
    .io_output(mac_15_30_io_output),
    .io_passthrough(mac_15_30_io_passthrough)
  );
  MAC mac_15_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_15_31_clock),
    .reset(mac_15_31_reset),
    .io_load(mac_15_31_io_load),
    .io_mulInput(mac_15_31_io_mulInput),
    .io_addInput(mac_15_31_io_addInput),
    .io_output(mac_15_31_io_output),
    .io_passthrough(mac_15_31_io_passthrough)
  );
  MAC mac_16_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_0_clock),
    .reset(mac_16_0_reset),
    .io_load(mac_16_0_io_load),
    .io_mulInput(mac_16_0_io_mulInput),
    .io_addInput(mac_16_0_io_addInput),
    .io_output(mac_16_0_io_output),
    .io_passthrough(mac_16_0_io_passthrough)
  );
  MAC mac_16_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_1_clock),
    .reset(mac_16_1_reset),
    .io_load(mac_16_1_io_load),
    .io_mulInput(mac_16_1_io_mulInput),
    .io_addInput(mac_16_1_io_addInput),
    .io_output(mac_16_1_io_output),
    .io_passthrough(mac_16_1_io_passthrough)
  );
  MAC mac_16_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_2_clock),
    .reset(mac_16_2_reset),
    .io_load(mac_16_2_io_load),
    .io_mulInput(mac_16_2_io_mulInput),
    .io_addInput(mac_16_2_io_addInput),
    .io_output(mac_16_2_io_output),
    .io_passthrough(mac_16_2_io_passthrough)
  );
  MAC mac_16_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_3_clock),
    .reset(mac_16_3_reset),
    .io_load(mac_16_3_io_load),
    .io_mulInput(mac_16_3_io_mulInput),
    .io_addInput(mac_16_3_io_addInput),
    .io_output(mac_16_3_io_output),
    .io_passthrough(mac_16_3_io_passthrough)
  );
  MAC mac_16_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_4_clock),
    .reset(mac_16_4_reset),
    .io_load(mac_16_4_io_load),
    .io_mulInput(mac_16_4_io_mulInput),
    .io_addInput(mac_16_4_io_addInput),
    .io_output(mac_16_4_io_output),
    .io_passthrough(mac_16_4_io_passthrough)
  );
  MAC mac_16_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_5_clock),
    .reset(mac_16_5_reset),
    .io_load(mac_16_5_io_load),
    .io_mulInput(mac_16_5_io_mulInput),
    .io_addInput(mac_16_5_io_addInput),
    .io_output(mac_16_5_io_output),
    .io_passthrough(mac_16_5_io_passthrough)
  );
  MAC mac_16_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_6_clock),
    .reset(mac_16_6_reset),
    .io_load(mac_16_6_io_load),
    .io_mulInput(mac_16_6_io_mulInput),
    .io_addInput(mac_16_6_io_addInput),
    .io_output(mac_16_6_io_output),
    .io_passthrough(mac_16_6_io_passthrough)
  );
  MAC mac_16_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_7_clock),
    .reset(mac_16_7_reset),
    .io_load(mac_16_7_io_load),
    .io_mulInput(mac_16_7_io_mulInput),
    .io_addInput(mac_16_7_io_addInput),
    .io_output(mac_16_7_io_output),
    .io_passthrough(mac_16_7_io_passthrough)
  );
  MAC mac_16_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_8_clock),
    .reset(mac_16_8_reset),
    .io_load(mac_16_8_io_load),
    .io_mulInput(mac_16_8_io_mulInput),
    .io_addInput(mac_16_8_io_addInput),
    .io_output(mac_16_8_io_output),
    .io_passthrough(mac_16_8_io_passthrough)
  );
  MAC mac_16_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_9_clock),
    .reset(mac_16_9_reset),
    .io_load(mac_16_9_io_load),
    .io_mulInput(mac_16_9_io_mulInput),
    .io_addInput(mac_16_9_io_addInput),
    .io_output(mac_16_9_io_output),
    .io_passthrough(mac_16_9_io_passthrough)
  );
  MAC mac_16_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_10_clock),
    .reset(mac_16_10_reset),
    .io_load(mac_16_10_io_load),
    .io_mulInput(mac_16_10_io_mulInput),
    .io_addInput(mac_16_10_io_addInput),
    .io_output(mac_16_10_io_output),
    .io_passthrough(mac_16_10_io_passthrough)
  );
  MAC mac_16_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_11_clock),
    .reset(mac_16_11_reset),
    .io_load(mac_16_11_io_load),
    .io_mulInput(mac_16_11_io_mulInput),
    .io_addInput(mac_16_11_io_addInput),
    .io_output(mac_16_11_io_output),
    .io_passthrough(mac_16_11_io_passthrough)
  );
  MAC mac_16_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_12_clock),
    .reset(mac_16_12_reset),
    .io_load(mac_16_12_io_load),
    .io_mulInput(mac_16_12_io_mulInput),
    .io_addInput(mac_16_12_io_addInput),
    .io_output(mac_16_12_io_output),
    .io_passthrough(mac_16_12_io_passthrough)
  );
  MAC mac_16_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_13_clock),
    .reset(mac_16_13_reset),
    .io_load(mac_16_13_io_load),
    .io_mulInput(mac_16_13_io_mulInput),
    .io_addInput(mac_16_13_io_addInput),
    .io_output(mac_16_13_io_output),
    .io_passthrough(mac_16_13_io_passthrough)
  );
  MAC mac_16_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_14_clock),
    .reset(mac_16_14_reset),
    .io_load(mac_16_14_io_load),
    .io_mulInput(mac_16_14_io_mulInput),
    .io_addInput(mac_16_14_io_addInput),
    .io_output(mac_16_14_io_output),
    .io_passthrough(mac_16_14_io_passthrough)
  );
  MAC mac_16_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_15_clock),
    .reset(mac_16_15_reset),
    .io_load(mac_16_15_io_load),
    .io_mulInput(mac_16_15_io_mulInput),
    .io_addInput(mac_16_15_io_addInput),
    .io_output(mac_16_15_io_output),
    .io_passthrough(mac_16_15_io_passthrough)
  );
  MAC mac_16_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_16_clock),
    .reset(mac_16_16_reset),
    .io_load(mac_16_16_io_load),
    .io_mulInput(mac_16_16_io_mulInput),
    .io_addInput(mac_16_16_io_addInput),
    .io_output(mac_16_16_io_output),
    .io_passthrough(mac_16_16_io_passthrough)
  );
  MAC mac_16_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_17_clock),
    .reset(mac_16_17_reset),
    .io_load(mac_16_17_io_load),
    .io_mulInput(mac_16_17_io_mulInput),
    .io_addInput(mac_16_17_io_addInput),
    .io_output(mac_16_17_io_output),
    .io_passthrough(mac_16_17_io_passthrough)
  );
  MAC mac_16_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_18_clock),
    .reset(mac_16_18_reset),
    .io_load(mac_16_18_io_load),
    .io_mulInput(mac_16_18_io_mulInput),
    .io_addInput(mac_16_18_io_addInput),
    .io_output(mac_16_18_io_output),
    .io_passthrough(mac_16_18_io_passthrough)
  );
  MAC mac_16_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_19_clock),
    .reset(mac_16_19_reset),
    .io_load(mac_16_19_io_load),
    .io_mulInput(mac_16_19_io_mulInput),
    .io_addInput(mac_16_19_io_addInput),
    .io_output(mac_16_19_io_output),
    .io_passthrough(mac_16_19_io_passthrough)
  );
  MAC mac_16_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_20_clock),
    .reset(mac_16_20_reset),
    .io_load(mac_16_20_io_load),
    .io_mulInput(mac_16_20_io_mulInput),
    .io_addInput(mac_16_20_io_addInput),
    .io_output(mac_16_20_io_output),
    .io_passthrough(mac_16_20_io_passthrough)
  );
  MAC mac_16_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_21_clock),
    .reset(mac_16_21_reset),
    .io_load(mac_16_21_io_load),
    .io_mulInput(mac_16_21_io_mulInput),
    .io_addInput(mac_16_21_io_addInput),
    .io_output(mac_16_21_io_output),
    .io_passthrough(mac_16_21_io_passthrough)
  );
  MAC mac_16_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_22_clock),
    .reset(mac_16_22_reset),
    .io_load(mac_16_22_io_load),
    .io_mulInput(mac_16_22_io_mulInput),
    .io_addInput(mac_16_22_io_addInput),
    .io_output(mac_16_22_io_output),
    .io_passthrough(mac_16_22_io_passthrough)
  );
  MAC mac_16_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_23_clock),
    .reset(mac_16_23_reset),
    .io_load(mac_16_23_io_load),
    .io_mulInput(mac_16_23_io_mulInput),
    .io_addInput(mac_16_23_io_addInput),
    .io_output(mac_16_23_io_output),
    .io_passthrough(mac_16_23_io_passthrough)
  );
  MAC mac_16_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_24_clock),
    .reset(mac_16_24_reset),
    .io_load(mac_16_24_io_load),
    .io_mulInput(mac_16_24_io_mulInput),
    .io_addInput(mac_16_24_io_addInput),
    .io_output(mac_16_24_io_output),
    .io_passthrough(mac_16_24_io_passthrough)
  );
  MAC mac_16_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_25_clock),
    .reset(mac_16_25_reset),
    .io_load(mac_16_25_io_load),
    .io_mulInput(mac_16_25_io_mulInput),
    .io_addInput(mac_16_25_io_addInput),
    .io_output(mac_16_25_io_output),
    .io_passthrough(mac_16_25_io_passthrough)
  );
  MAC mac_16_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_26_clock),
    .reset(mac_16_26_reset),
    .io_load(mac_16_26_io_load),
    .io_mulInput(mac_16_26_io_mulInput),
    .io_addInput(mac_16_26_io_addInput),
    .io_output(mac_16_26_io_output),
    .io_passthrough(mac_16_26_io_passthrough)
  );
  MAC mac_16_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_27_clock),
    .reset(mac_16_27_reset),
    .io_load(mac_16_27_io_load),
    .io_mulInput(mac_16_27_io_mulInput),
    .io_addInput(mac_16_27_io_addInput),
    .io_output(mac_16_27_io_output),
    .io_passthrough(mac_16_27_io_passthrough)
  );
  MAC mac_16_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_28_clock),
    .reset(mac_16_28_reset),
    .io_load(mac_16_28_io_load),
    .io_mulInput(mac_16_28_io_mulInput),
    .io_addInput(mac_16_28_io_addInput),
    .io_output(mac_16_28_io_output),
    .io_passthrough(mac_16_28_io_passthrough)
  );
  MAC mac_16_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_29_clock),
    .reset(mac_16_29_reset),
    .io_load(mac_16_29_io_load),
    .io_mulInput(mac_16_29_io_mulInput),
    .io_addInput(mac_16_29_io_addInput),
    .io_output(mac_16_29_io_output),
    .io_passthrough(mac_16_29_io_passthrough)
  );
  MAC mac_16_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_30_clock),
    .reset(mac_16_30_reset),
    .io_load(mac_16_30_io_load),
    .io_mulInput(mac_16_30_io_mulInput),
    .io_addInput(mac_16_30_io_addInput),
    .io_output(mac_16_30_io_output),
    .io_passthrough(mac_16_30_io_passthrough)
  );
  MAC mac_16_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_16_31_clock),
    .reset(mac_16_31_reset),
    .io_load(mac_16_31_io_load),
    .io_mulInput(mac_16_31_io_mulInput),
    .io_addInput(mac_16_31_io_addInput),
    .io_output(mac_16_31_io_output),
    .io_passthrough(mac_16_31_io_passthrough)
  );
  MAC mac_17_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_0_clock),
    .reset(mac_17_0_reset),
    .io_load(mac_17_0_io_load),
    .io_mulInput(mac_17_0_io_mulInput),
    .io_addInput(mac_17_0_io_addInput),
    .io_output(mac_17_0_io_output),
    .io_passthrough(mac_17_0_io_passthrough)
  );
  MAC mac_17_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_1_clock),
    .reset(mac_17_1_reset),
    .io_load(mac_17_1_io_load),
    .io_mulInput(mac_17_1_io_mulInput),
    .io_addInput(mac_17_1_io_addInput),
    .io_output(mac_17_1_io_output),
    .io_passthrough(mac_17_1_io_passthrough)
  );
  MAC mac_17_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_2_clock),
    .reset(mac_17_2_reset),
    .io_load(mac_17_2_io_load),
    .io_mulInput(mac_17_2_io_mulInput),
    .io_addInput(mac_17_2_io_addInput),
    .io_output(mac_17_2_io_output),
    .io_passthrough(mac_17_2_io_passthrough)
  );
  MAC mac_17_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_3_clock),
    .reset(mac_17_3_reset),
    .io_load(mac_17_3_io_load),
    .io_mulInput(mac_17_3_io_mulInput),
    .io_addInput(mac_17_3_io_addInput),
    .io_output(mac_17_3_io_output),
    .io_passthrough(mac_17_3_io_passthrough)
  );
  MAC mac_17_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_4_clock),
    .reset(mac_17_4_reset),
    .io_load(mac_17_4_io_load),
    .io_mulInput(mac_17_4_io_mulInput),
    .io_addInput(mac_17_4_io_addInput),
    .io_output(mac_17_4_io_output),
    .io_passthrough(mac_17_4_io_passthrough)
  );
  MAC mac_17_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_5_clock),
    .reset(mac_17_5_reset),
    .io_load(mac_17_5_io_load),
    .io_mulInput(mac_17_5_io_mulInput),
    .io_addInput(mac_17_5_io_addInput),
    .io_output(mac_17_5_io_output),
    .io_passthrough(mac_17_5_io_passthrough)
  );
  MAC mac_17_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_6_clock),
    .reset(mac_17_6_reset),
    .io_load(mac_17_6_io_load),
    .io_mulInput(mac_17_6_io_mulInput),
    .io_addInput(mac_17_6_io_addInput),
    .io_output(mac_17_6_io_output),
    .io_passthrough(mac_17_6_io_passthrough)
  );
  MAC mac_17_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_7_clock),
    .reset(mac_17_7_reset),
    .io_load(mac_17_7_io_load),
    .io_mulInput(mac_17_7_io_mulInput),
    .io_addInput(mac_17_7_io_addInput),
    .io_output(mac_17_7_io_output),
    .io_passthrough(mac_17_7_io_passthrough)
  );
  MAC mac_17_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_8_clock),
    .reset(mac_17_8_reset),
    .io_load(mac_17_8_io_load),
    .io_mulInput(mac_17_8_io_mulInput),
    .io_addInput(mac_17_8_io_addInput),
    .io_output(mac_17_8_io_output),
    .io_passthrough(mac_17_8_io_passthrough)
  );
  MAC mac_17_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_9_clock),
    .reset(mac_17_9_reset),
    .io_load(mac_17_9_io_load),
    .io_mulInput(mac_17_9_io_mulInput),
    .io_addInput(mac_17_9_io_addInput),
    .io_output(mac_17_9_io_output),
    .io_passthrough(mac_17_9_io_passthrough)
  );
  MAC mac_17_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_10_clock),
    .reset(mac_17_10_reset),
    .io_load(mac_17_10_io_load),
    .io_mulInput(mac_17_10_io_mulInput),
    .io_addInput(mac_17_10_io_addInput),
    .io_output(mac_17_10_io_output),
    .io_passthrough(mac_17_10_io_passthrough)
  );
  MAC mac_17_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_11_clock),
    .reset(mac_17_11_reset),
    .io_load(mac_17_11_io_load),
    .io_mulInput(mac_17_11_io_mulInput),
    .io_addInput(mac_17_11_io_addInput),
    .io_output(mac_17_11_io_output),
    .io_passthrough(mac_17_11_io_passthrough)
  );
  MAC mac_17_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_12_clock),
    .reset(mac_17_12_reset),
    .io_load(mac_17_12_io_load),
    .io_mulInput(mac_17_12_io_mulInput),
    .io_addInput(mac_17_12_io_addInput),
    .io_output(mac_17_12_io_output),
    .io_passthrough(mac_17_12_io_passthrough)
  );
  MAC mac_17_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_13_clock),
    .reset(mac_17_13_reset),
    .io_load(mac_17_13_io_load),
    .io_mulInput(mac_17_13_io_mulInput),
    .io_addInput(mac_17_13_io_addInput),
    .io_output(mac_17_13_io_output),
    .io_passthrough(mac_17_13_io_passthrough)
  );
  MAC mac_17_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_14_clock),
    .reset(mac_17_14_reset),
    .io_load(mac_17_14_io_load),
    .io_mulInput(mac_17_14_io_mulInput),
    .io_addInput(mac_17_14_io_addInput),
    .io_output(mac_17_14_io_output),
    .io_passthrough(mac_17_14_io_passthrough)
  );
  MAC mac_17_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_15_clock),
    .reset(mac_17_15_reset),
    .io_load(mac_17_15_io_load),
    .io_mulInput(mac_17_15_io_mulInput),
    .io_addInput(mac_17_15_io_addInput),
    .io_output(mac_17_15_io_output),
    .io_passthrough(mac_17_15_io_passthrough)
  );
  MAC mac_17_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_16_clock),
    .reset(mac_17_16_reset),
    .io_load(mac_17_16_io_load),
    .io_mulInput(mac_17_16_io_mulInput),
    .io_addInput(mac_17_16_io_addInput),
    .io_output(mac_17_16_io_output),
    .io_passthrough(mac_17_16_io_passthrough)
  );
  MAC mac_17_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_17_clock),
    .reset(mac_17_17_reset),
    .io_load(mac_17_17_io_load),
    .io_mulInput(mac_17_17_io_mulInput),
    .io_addInput(mac_17_17_io_addInput),
    .io_output(mac_17_17_io_output),
    .io_passthrough(mac_17_17_io_passthrough)
  );
  MAC mac_17_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_18_clock),
    .reset(mac_17_18_reset),
    .io_load(mac_17_18_io_load),
    .io_mulInput(mac_17_18_io_mulInput),
    .io_addInput(mac_17_18_io_addInput),
    .io_output(mac_17_18_io_output),
    .io_passthrough(mac_17_18_io_passthrough)
  );
  MAC mac_17_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_19_clock),
    .reset(mac_17_19_reset),
    .io_load(mac_17_19_io_load),
    .io_mulInput(mac_17_19_io_mulInput),
    .io_addInput(mac_17_19_io_addInput),
    .io_output(mac_17_19_io_output),
    .io_passthrough(mac_17_19_io_passthrough)
  );
  MAC mac_17_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_20_clock),
    .reset(mac_17_20_reset),
    .io_load(mac_17_20_io_load),
    .io_mulInput(mac_17_20_io_mulInput),
    .io_addInput(mac_17_20_io_addInput),
    .io_output(mac_17_20_io_output),
    .io_passthrough(mac_17_20_io_passthrough)
  );
  MAC mac_17_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_21_clock),
    .reset(mac_17_21_reset),
    .io_load(mac_17_21_io_load),
    .io_mulInput(mac_17_21_io_mulInput),
    .io_addInput(mac_17_21_io_addInput),
    .io_output(mac_17_21_io_output),
    .io_passthrough(mac_17_21_io_passthrough)
  );
  MAC mac_17_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_22_clock),
    .reset(mac_17_22_reset),
    .io_load(mac_17_22_io_load),
    .io_mulInput(mac_17_22_io_mulInput),
    .io_addInput(mac_17_22_io_addInput),
    .io_output(mac_17_22_io_output),
    .io_passthrough(mac_17_22_io_passthrough)
  );
  MAC mac_17_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_23_clock),
    .reset(mac_17_23_reset),
    .io_load(mac_17_23_io_load),
    .io_mulInput(mac_17_23_io_mulInput),
    .io_addInput(mac_17_23_io_addInput),
    .io_output(mac_17_23_io_output),
    .io_passthrough(mac_17_23_io_passthrough)
  );
  MAC mac_17_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_24_clock),
    .reset(mac_17_24_reset),
    .io_load(mac_17_24_io_load),
    .io_mulInput(mac_17_24_io_mulInput),
    .io_addInput(mac_17_24_io_addInput),
    .io_output(mac_17_24_io_output),
    .io_passthrough(mac_17_24_io_passthrough)
  );
  MAC mac_17_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_25_clock),
    .reset(mac_17_25_reset),
    .io_load(mac_17_25_io_load),
    .io_mulInput(mac_17_25_io_mulInput),
    .io_addInput(mac_17_25_io_addInput),
    .io_output(mac_17_25_io_output),
    .io_passthrough(mac_17_25_io_passthrough)
  );
  MAC mac_17_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_26_clock),
    .reset(mac_17_26_reset),
    .io_load(mac_17_26_io_load),
    .io_mulInput(mac_17_26_io_mulInput),
    .io_addInput(mac_17_26_io_addInput),
    .io_output(mac_17_26_io_output),
    .io_passthrough(mac_17_26_io_passthrough)
  );
  MAC mac_17_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_27_clock),
    .reset(mac_17_27_reset),
    .io_load(mac_17_27_io_load),
    .io_mulInput(mac_17_27_io_mulInput),
    .io_addInput(mac_17_27_io_addInput),
    .io_output(mac_17_27_io_output),
    .io_passthrough(mac_17_27_io_passthrough)
  );
  MAC mac_17_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_28_clock),
    .reset(mac_17_28_reset),
    .io_load(mac_17_28_io_load),
    .io_mulInput(mac_17_28_io_mulInput),
    .io_addInput(mac_17_28_io_addInput),
    .io_output(mac_17_28_io_output),
    .io_passthrough(mac_17_28_io_passthrough)
  );
  MAC mac_17_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_29_clock),
    .reset(mac_17_29_reset),
    .io_load(mac_17_29_io_load),
    .io_mulInput(mac_17_29_io_mulInput),
    .io_addInput(mac_17_29_io_addInput),
    .io_output(mac_17_29_io_output),
    .io_passthrough(mac_17_29_io_passthrough)
  );
  MAC mac_17_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_30_clock),
    .reset(mac_17_30_reset),
    .io_load(mac_17_30_io_load),
    .io_mulInput(mac_17_30_io_mulInput),
    .io_addInput(mac_17_30_io_addInput),
    .io_output(mac_17_30_io_output),
    .io_passthrough(mac_17_30_io_passthrough)
  );
  MAC mac_17_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_17_31_clock),
    .reset(mac_17_31_reset),
    .io_load(mac_17_31_io_load),
    .io_mulInput(mac_17_31_io_mulInput),
    .io_addInput(mac_17_31_io_addInput),
    .io_output(mac_17_31_io_output),
    .io_passthrough(mac_17_31_io_passthrough)
  );
  MAC mac_18_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_0_clock),
    .reset(mac_18_0_reset),
    .io_load(mac_18_0_io_load),
    .io_mulInput(mac_18_0_io_mulInput),
    .io_addInput(mac_18_0_io_addInput),
    .io_output(mac_18_0_io_output),
    .io_passthrough(mac_18_0_io_passthrough)
  );
  MAC mac_18_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_1_clock),
    .reset(mac_18_1_reset),
    .io_load(mac_18_1_io_load),
    .io_mulInput(mac_18_1_io_mulInput),
    .io_addInput(mac_18_1_io_addInput),
    .io_output(mac_18_1_io_output),
    .io_passthrough(mac_18_1_io_passthrough)
  );
  MAC mac_18_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_2_clock),
    .reset(mac_18_2_reset),
    .io_load(mac_18_2_io_load),
    .io_mulInput(mac_18_2_io_mulInput),
    .io_addInput(mac_18_2_io_addInput),
    .io_output(mac_18_2_io_output),
    .io_passthrough(mac_18_2_io_passthrough)
  );
  MAC mac_18_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_3_clock),
    .reset(mac_18_3_reset),
    .io_load(mac_18_3_io_load),
    .io_mulInput(mac_18_3_io_mulInput),
    .io_addInput(mac_18_3_io_addInput),
    .io_output(mac_18_3_io_output),
    .io_passthrough(mac_18_3_io_passthrough)
  );
  MAC mac_18_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_4_clock),
    .reset(mac_18_4_reset),
    .io_load(mac_18_4_io_load),
    .io_mulInput(mac_18_4_io_mulInput),
    .io_addInput(mac_18_4_io_addInput),
    .io_output(mac_18_4_io_output),
    .io_passthrough(mac_18_4_io_passthrough)
  );
  MAC mac_18_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_5_clock),
    .reset(mac_18_5_reset),
    .io_load(mac_18_5_io_load),
    .io_mulInput(mac_18_5_io_mulInput),
    .io_addInput(mac_18_5_io_addInput),
    .io_output(mac_18_5_io_output),
    .io_passthrough(mac_18_5_io_passthrough)
  );
  MAC mac_18_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_6_clock),
    .reset(mac_18_6_reset),
    .io_load(mac_18_6_io_load),
    .io_mulInput(mac_18_6_io_mulInput),
    .io_addInput(mac_18_6_io_addInput),
    .io_output(mac_18_6_io_output),
    .io_passthrough(mac_18_6_io_passthrough)
  );
  MAC mac_18_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_7_clock),
    .reset(mac_18_7_reset),
    .io_load(mac_18_7_io_load),
    .io_mulInput(mac_18_7_io_mulInput),
    .io_addInput(mac_18_7_io_addInput),
    .io_output(mac_18_7_io_output),
    .io_passthrough(mac_18_7_io_passthrough)
  );
  MAC mac_18_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_8_clock),
    .reset(mac_18_8_reset),
    .io_load(mac_18_8_io_load),
    .io_mulInput(mac_18_8_io_mulInput),
    .io_addInput(mac_18_8_io_addInput),
    .io_output(mac_18_8_io_output),
    .io_passthrough(mac_18_8_io_passthrough)
  );
  MAC mac_18_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_9_clock),
    .reset(mac_18_9_reset),
    .io_load(mac_18_9_io_load),
    .io_mulInput(mac_18_9_io_mulInput),
    .io_addInput(mac_18_9_io_addInput),
    .io_output(mac_18_9_io_output),
    .io_passthrough(mac_18_9_io_passthrough)
  );
  MAC mac_18_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_10_clock),
    .reset(mac_18_10_reset),
    .io_load(mac_18_10_io_load),
    .io_mulInput(mac_18_10_io_mulInput),
    .io_addInput(mac_18_10_io_addInput),
    .io_output(mac_18_10_io_output),
    .io_passthrough(mac_18_10_io_passthrough)
  );
  MAC mac_18_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_11_clock),
    .reset(mac_18_11_reset),
    .io_load(mac_18_11_io_load),
    .io_mulInput(mac_18_11_io_mulInput),
    .io_addInput(mac_18_11_io_addInput),
    .io_output(mac_18_11_io_output),
    .io_passthrough(mac_18_11_io_passthrough)
  );
  MAC mac_18_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_12_clock),
    .reset(mac_18_12_reset),
    .io_load(mac_18_12_io_load),
    .io_mulInput(mac_18_12_io_mulInput),
    .io_addInput(mac_18_12_io_addInput),
    .io_output(mac_18_12_io_output),
    .io_passthrough(mac_18_12_io_passthrough)
  );
  MAC mac_18_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_13_clock),
    .reset(mac_18_13_reset),
    .io_load(mac_18_13_io_load),
    .io_mulInput(mac_18_13_io_mulInput),
    .io_addInput(mac_18_13_io_addInput),
    .io_output(mac_18_13_io_output),
    .io_passthrough(mac_18_13_io_passthrough)
  );
  MAC mac_18_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_14_clock),
    .reset(mac_18_14_reset),
    .io_load(mac_18_14_io_load),
    .io_mulInput(mac_18_14_io_mulInput),
    .io_addInput(mac_18_14_io_addInput),
    .io_output(mac_18_14_io_output),
    .io_passthrough(mac_18_14_io_passthrough)
  );
  MAC mac_18_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_15_clock),
    .reset(mac_18_15_reset),
    .io_load(mac_18_15_io_load),
    .io_mulInput(mac_18_15_io_mulInput),
    .io_addInput(mac_18_15_io_addInput),
    .io_output(mac_18_15_io_output),
    .io_passthrough(mac_18_15_io_passthrough)
  );
  MAC mac_18_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_16_clock),
    .reset(mac_18_16_reset),
    .io_load(mac_18_16_io_load),
    .io_mulInput(mac_18_16_io_mulInput),
    .io_addInput(mac_18_16_io_addInput),
    .io_output(mac_18_16_io_output),
    .io_passthrough(mac_18_16_io_passthrough)
  );
  MAC mac_18_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_17_clock),
    .reset(mac_18_17_reset),
    .io_load(mac_18_17_io_load),
    .io_mulInput(mac_18_17_io_mulInput),
    .io_addInput(mac_18_17_io_addInput),
    .io_output(mac_18_17_io_output),
    .io_passthrough(mac_18_17_io_passthrough)
  );
  MAC mac_18_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_18_clock),
    .reset(mac_18_18_reset),
    .io_load(mac_18_18_io_load),
    .io_mulInput(mac_18_18_io_mulInput),
    .io_addInput(mac_18_18_io_addInput),
    .io_output(mac_18_18_io_output),
    .io_passthrough(mac_18_18_io_passthrough)
  );
  MAC mac_18_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_19_clock),
    .reset(mac_18_19_reset),
    .io_load(mac_18_19_io_load),
    .io_mulInput(mac_18_19_io_mulInput),
    .io_addInput(mac_18_19_io_addInput),
    .io_output(mac_18_19_io_output),
    .io_passthrough(mac_18_19_io_passthrough)
  );
  MAC mac_18_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_20_clock),
    .reset(mac_18_20_reset),
    .io_load(mac_18_20_io_load),
    .io_mulInput(mac_18_20_io_mulInput),
    .io_addInput(mac_18_20_io_addInput),
    .io_output(mac_18_20_io_output),
    .io_passthrough(mac_18_20_io_passthrough)
  );
  MAC mac_18_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_21_clock),
    .reset(mac_18_21_reset),
    .io_load(mac_18_21_io_load),
    .io_mulInput(mac_18_21_io_mulInput),
    .io_addInput(mac_18_21_io_addInput),
    .io_output(mac_18_21_io_output),
    .io_passthrough(mac_18_21_io_passthrough)
  );
  MAC mac_18_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_22_clock),
    .reset(mac_18_22_reset),
    .io_load(mac_18_22_io_load),
    .io_mulInput(mac_18_22_io_mulInput),
    .io_addInput(mac_18_22_io_addInput),
    .io_output(mac_18_22_io_output),
    .io_passthrough(mac_18_22_io_passthrough)
  );
  MAC mac_18_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_23_clock),
    .reset(mac_18_23_reset),
    .io_load(mac_18_23_io_load),
    .io_mulInput(mac_18_23_io_mulInput),
    .io_addInput(mac_18_23_io_addInput),
    .io_output(mac_18_23_io_output),
    .io_passthrough(mac_18_23_io_passthrough)
  );
  MAC mac_18_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_24_clock),
    .reset(mac_18_24_reset),
    .io_load(mac_18_24_io_load),
    .io_mulInput(mac_18_24_io_mulInput),
    .io_addInput(mac_18_24_io_addInput),
    .io_output(mac_18_24_io_output),
    .io_passthrough(mac_18_24_io_passthrough)
  );
  MAC mac_18_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_25_clock),
    .reset(mac_18_25_reset),
    .io_load(mac_18_25_io_load),
    .io_mulInput(mac_18_25_io_mulInput),
    .io_addInput(mac_18_25_io_addInput),
    .io_output(mac_18_25_io_output),
    .io_passthrough(mac_18_25_io_passthrough)
  );
  MAC mac_18_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_26_clock),
    .reset(mac_18_26_reset),
    .io_load(mac_18_26_io_load),
    .io_mulInput(mac_18_26_io_mulInput),
    .io_addInput(mac_18_26_io_addInput),
    .io_output(mac_18_26_io_output),
    .io_passthrough(mac_18_26_io_passthrough)
  );
  MAC mac_18_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_27_clock),
    .reset(mac_18_27_reset),
    .io_load(mac_18_27_io_load),
    .io_mulInput(mac_18_27_io_mulInput),
    .io_addInput(mac_18_27_io_addInput),
    .io_output(mac_18_27_io_output),
    .io_passthrough(mac_18_27_io_passthrough)
  );
  MAC mac_18_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_28_clock),
    .reset(mac_18_28_reset),
    .io_load(mac_18_28_io_load),
    .io_mulInput(mac_18_28_io_mulInput),
    .io_addInput(mac_18_28_io_addInput),
    .io_output(mac_18_28_io_output),
    .io_passthrough(mac_18_28_io_passthrough)
  );
  MAC mac_18_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_29_clock),
    .reset(mac_18_29_reset),
    .io_load(mac_18_29_io_load),
    .io_mulInput(mac_18_29_io_mulInput),
    .io_addInput(mac_18_29_io_addInput),
    .io_output(mac_18_29_io_output),
    .io_passthrough(mac_18_29_io_passthrough)
  );
  MAC mac_18_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_30_clock),
    .reset(mac_18_30_reset),
    .io_load(mac_18_30_io_load),
    .io_mulInput(mac_18_30_io_mulInput),
    .io_addInput(mac_18_30_io_addInput),
    .io_output(mac_18_30_io_output),
    .io_passthrough(mac_18_30_io_passthrough)
  );
  MAC mac_18_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_18_31_clock),
    .reset(mac_18_31_reset),
    .io_load(mac_18_31_io_load),
    .io_mulInput(mac_18_31_io_mulInput),
    .io_addInput(mac_18_31_io_addInput),
    .io_output(mac_18_31_io_output),
    .io_passthrough(mac_18_31_io_passthrough)
  );
  MAC mac_19_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_0_clock),
    .reset(mac_19_0_reset),
    .io_load(mac_19_0_io_load),
    .io_mulInput(mac_19_0_io_mulInput),
    .io_addInput(mac_19_0_io_addInput),
    .io_output(mac_19_0_io_output),
    .io_passthrough(mac_19_0_io_passthrough)
  );
  MAC mac_19_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_1_clock),
    .reset(mac_19_1_reset),
    .io_load(mac_19_1_io_load),
    .io_mulInput(mac_19_1_io_mulInput),
    .io_addInput(mac_19_1_io_addInput),
    .io_output(mac_19_1_io_output),
    .io_passthrough(mac_19_1_io_passthrough)
  );
  MAC mac_19_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_2_clock),
    .reset(mac_19_2_reset),
    .io_load(mac_19_2_io_load),
    .io_mulInput(mac_19_2_io_mulInput),
    .io_addInput(mac_19_2_io_addInput),
    .io_output(mac_19_2_io_output),
    .io_passthrough(mac_19_2_io_passthrough)
  );
  MAC mac_19_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_3_clock),
    .reset(mac_19_3_reset),
    .io_load(mac_19_3_io_load),
    .io_mulInput(mac_19_3_io_mulInput),
    .io_addInput(mac_19_3_io_addInput),
    .io_output(mac_19_3_io_output),
    .io_passthrough(mac_19_3_io_passthrough)
  );
  MAC mac_19_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_4_clock),
    .reset(mac_19_4_reset),
    .io_load(mac_19_4_io_load),
    .io_mulInput(mac_19_4_io_mulInput),
    .io_addInput(mac_19_4_io_addInput),
    .io_output(mac_19_4_io_output),
    .io_passthrough(mac_19_4_io_passthrough)
  );
  MAC mac_19_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_5_clock),
    .reset(mac_19_5_reset),
    .io_load(mac_19_5_io_load),
    .io_mulInput(mac_19_5_io_mulInput),
    .io_addInput(mac_19_5_io_addInput),
    .io_output(mac_19_5_io_output),
    .io_passthrough(mac_19_5_io_passthrough)
  );
  MAC mac_19_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_6_clock),
    .reset(mac_19_6_reset),
    .io_load(mac_19_6_io_load),
    .io_mulInput(mac_19_6_io_mulInput),
    .io_addInput(mac_19_6_io_addInput),
    .io_output(mac_19_6_io_output),
    .io_passthrough(mac_19_6_io_passthrough)
  );
  MAC mac_19_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_7_clock),
    .reset(mac_19_7_reset),
    .io_load(mac_19_7_io_load),
    .io_mulInput(mac_19_7_io_mulInput),
    .io_addInput(mac_19_7_io_addInput),
    .io_output(mac_19_7_io_output),
    .io_passthrough(mac_19_7_io_passthrough)
  );
  MAC mac_19_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_8_clock),
    .reset(mac_19_8_reset),
    .io_load(mac_19_8_io_load),
    .io_mulInput(mac_19_8_io_mulInput),
    .io_addInput(mac_19_8_io_addInput),
    .io_output(mac_19_8_io_output),
    .io_passthrough(mac_19_8_io_passthrough)
  );
  MAC mac_19_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_9_clock),
    .reset(mac_19_9_reset),
    .io_load(mac_19_9_io_load),
    .io_mulInput(mac_19_9_io_mulInput),
    .io_addInput(mac_19_9_io_addInput),
    .io_output(mac_19_9_io_output),
    .io_passthrough(mac_19_9_io_passthrough)
  );
  MAC mac_19_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_10_clock),
    .reset(mac_19_10_reset),
    .io_load(mac_19_10_io_load),
    .io_mulInput(mac_19_10_io_mulInput),
    .io_addInput(mac_19_10_io_addInput),
    .io_output(mac_19_10_io_output),
    .io_passthrough(mac_19_10_io_passthrough)
  );
  MAC mac_19_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_11_clock),
    .reset(mac_19_11_reset),
    .io_load(mac_19_11_io_load),
    .io_mulInput(mac_19_11_io_mulInput),
    .io_addInput(mac_19_11_io_addInput),
    .io_output(mac_19_11_io_output),
    .io_passthrough(mac_19_11_io_passthrough)
  );
  MAC mac_19_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_12_clock),
    .reset(mac_19_12_reset),
    .io_load(mac_19_12_io_load),
    .io_mulInput(mac_19_12_io_mulInput),
    .io_addInput(mac_19_12_io_addInput),
    .io_output(mac_19_12_io_output),
    .io_passthrough(mac_19_12_io_passthrough)
  );
  MAC mac_19_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_13_clock),
    .reset(mac_19_13_reset),
    .io_load(mac_19_13_io_load),
    .io_mulInput(mac_19_13_io_mulInput),
    .io_addInput(mac_19_13_io_addInput),
    .io_output(mac_19_13_io_output),
    .io_passthrough(mac_19_13_io_passthrough)
  );
  MAC mac_19_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_14_clock),
    .reset(mac_19_14_reset),
    .io_load(mac_19_14_io_load),
    .io_mulInput(mac_19_14_io_mulInput),
    .io_addInput(mac_19_14_io_addInput),
    .io_output(mac_19_14_io_output),
    .io_passthrough(mac_19_14_io_passthrough)
  );
  MAC mac_19_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_15_clock),
    .reset(mac_19_15_reset),
    .io_load(mac_19_15_io_load),
    .io_mulInput(mac_19_15_io_mulInput),
    .io_addInput(mac_19_15_io_addInput),
    .io_output(mac_19_15_io_output),
    .io_passthrough(mac_19_15_io_passthrough)
  );
  MAC mac_19_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_16_clock),
    .reset(mac_19_16_reset),
    .io_load(mac_19_16_io_load),
    .io_mulInput(mac_19_16_io_mulInput),
    .io_addInput(mac_19_16_io_addInput),
    .io_output(mac_19_16_io_output),
    .io_passthrough(mac_19_16_io_passthrough)
  );
  MAC mac_19_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_17_clock),
    .reset(mac_19_17_reset),
    .io_load(mac_19_17_io_load),
    .io_mulInput(mac_19_17_io_mulInput),
    .io_addInput(mac_19_17_io_addInput),
    .io_output(mac_19_17_io_output),
    .io_passthrough(mac_19_17_io_passthrough)
  );
  MAC mac_19_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_18_clock),
    .reset(mac_19_18_reset),
    .io_load(mac_19_18_io_load),
    .io_mulInput(mac_19_18_io_mulInput),
    .io_addInput(mac_19_18_io_addInput),
    .io_output(mac_19_18_io_output),
    .io_passthrough(mac_19_18_io_passthrough)
  );
  MAC mac_19_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_19_clock),
    .reset(mac_19_19_reset),
    .io_load(mac_19_19_io_load),
    .io_mulInput(mac_19_19_io_mulInput),
    .io_addInput(mac_19_19_io_addInput),
    .io_output(mac_19_19_io_output),
    .io_passthrough(mac_19_19_io_passthrough)
  );
  MAC mac_19_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_20_clock),
    .reset(mac_19_20_reset),
    .io_load(mac_19_20_io_load),
    .io_mulInput(mac_19_20_io_mulInput),
    .io_addInput(mac_19_20_io_addInput),
    .io_output(mac_19_20_io_output),
    .io_passthrough(mac_19_20_io_passthrough)
  );
  MAC mac_19_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_21_clock),
    .reset(mac_19_21_reset),
    .io_load(mac_19_21_io_load),
    .io_mulInput(mac_19_21_io_mulInput),
    .io_addInput(mac_19_21_io_addInput),
    .io_output(mac_19_21_io_output),
    .io_passthrough(mac_19_21_io_passthrough)
  );
  MAC mac_19_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_22_clock),
    .reset(mac_19_22_reset),
    .io_load(mac_19_22_io_load),
    .io_mulInput(mac_19_22_io_mulInput),
    .io_addInput(mac_19_22_io_addInput),
    .io_output(mac_19_22_io_output),
    .io_passthrough(mac_19_22_io_passthrough)
  );
  MAC mac_19_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_23_clock),
    .reset(mac_19_23_reset),
    .io_load(mac_19_23_io_load),
    .io_mulInput(mac_19_23_io_mulInput),
    .io_addInput(mac_19_23_io_addInput),
    .io_output(mac_19_23_io_output),
    .io_passthrough(mac_19_23_io_passthrough)
  );
  MAC mac_19_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_24_clock),
    .reset(mac_19_24_reset),
    .io_load(mac_19_24_io_load),
    .io_mulInput(mac_19_24_io_mulInput),
    .io_addInput(mac_19_24_io_addInput),
    .io_output(mac_19_24_io_output),
    .io_passthrough(mac_19_24_io_passthrough)
  );
  MAC mac_19_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_25_clock),
    .reset(mac_19_25_reset),
    .io_load(mac_19_25_io_load),
    .io_mulInput(mac_19_25_io_mulInput),
    .io_addInput(mac_19_25_io_addInput),
    .io_output(mac_19_25_io_output),
    .io_passthrough(mac_19_25_io_passthrough)
  );
  MAC mac_19_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_26_clock),
    .reset(mac_19_26_reset),
    .io_load(mac_19_26_io_load),
    .io_mulInput(mac_19_26_io_mulInput),
    .io_addInput(mac_19_26_io_addInput),
    .io_output(mac_19_26_io_output),
    .io_passthrough(mac_19_26_io_passthrough)
  );
  MAC mac_19_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_27_clock),
    .reset(mac_19_27_reset),
    .io_load(mac_19_27_io_load),
    .io_mulInput(mac_19_27_io_mulInput),
    .io_addInput(mac_19_27_io_addInput),
    .io_output(mac_19_27_io_output),
    .io_passthrough(mac_19_27_io_passthrough)
  );
  MAC mac_19_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_28_clock),
    .reset(mac_19_28_reset),
    .io_load(mac_19_28_io_load),
    .io_mulInput(mac_19_28_io_mulInput),
    .io_addInput(mac_19_28_io_addInput),
    .io_output(mac_19_28_io_output),
    .io_passthrough(mac_19_28_io_passthrough)
  );
  MAC mac_19_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_29_clock),
    .reset(mac_19_29_reset),
    .io_load(mac_19_29_io_load),
    .io_mulInput(mac_19_29_io_mulInput),
    .io_addInput(mac_19_29_io_addInput),
    .io_output(mac_19_29_io_output),
    .io_passthrough(mac_19_29_io_passthrough)
  );
  MAC mac_19_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_30_clock),
    .reset(mac_19_30_reset),
    .io_load(mac_19_30_io_load),
    .io_mulInput(mac_19_30_io_mulInput),
    .io_addInput(mac_19_30_io_addInput),
    .io_output(mac_19_30_io_output),
    .io_passthrough(mac_19_30_io_passthrough)
  );
  MAC mac_19_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_19_31_clock),
    .reset(mac_19_31_reset),
    .io_load(mac_19_31_io_load),
    .io_mulInput(mac_19_31_io_mulInput),
    .io_addInput(mac_19_31_io_addInput),
    .io_output(mac_19_31_io_output),
    .io_passthrough(mac_19_31_io_passthrough)
  );
  MAC mac_20_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_0_clock),
    .reset(mac_20_0_reset),
    .io_load(mac_20_0_io_load),
    .io_mulInput(mac_20_0_io_mulInput),
    .io_addInput(mac_20_0_io_addInput),
    .io_output(mac_20_0_io_output),
    .io_passthrough(mac_20_0_io_passthrough)
  );
  MAC mac_20_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_1_clock),
    .reset(mac_20_1_reset),
    .io_load(mac_20_1_io_load),
    .io_mulInput(mac_20_1_io_mulInput),
    .io_addInput(mac_20_1_io_addInput),
    .io_output(mac_20_1_io_output),
    .io_passthrough(mac_20_1_io_passthrough)
  );
  MAC mac_20_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_2_clock),
    .reset(mac_20_2_reset),
    .io_load(mac_20_2_io_load),
    .io_mulInput(mac_20_2_io_mulInput),
    .io_addInput(mac_20_2_io_addInput),
    .io_output(mac_20_2_io_output),
    .io_passthrough(mac_20_2_io_passthrough)
  );
  MAC mac_20_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_3_clock),
    .reset(mac_20_3_reset),
    .io_load(mac_20_3_io_load),
    .io_mulInput(mac_20_3_io_mulInput),
    .io_addInput(mac_20_3_io_addInput),
    .io_output(mac_20_3_io_output),
    .io_passthrough(mac_20_3_io_passthrough)
  );
  MAC mac_20_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_4_clock),
    .reset(mac_20_4_reset),
    .io_load(mac_20_4_io_load),
    .io_mulInput(mac_20_4_io_mulInput),
    .io_addInput(mac_20_4_io_addInput),
    .io_output(mac_20_4_io_output),
    .io_passthrough(mac_20_4_io_passthrough)
  );
  MAC mac_20_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_5_clock),
    .reset(mac_20_5_reset),
    .io_load(mac_20_5_io_load),
    .io_mulInput(mac_20_5_io_mulInput),
    .io_addInput(mac_20_5_io_addInput),
    .io_output(mac_20_5_io_output),
    .io_passthrough(mac_20_5_io_passthrough)
  );
  MAC mac_20_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_6_clock),
    .reset(mac_20_6_reset),
    .io_load(mac_20_6_io_load),
    .io_mulInput(mac_20_6_io_mulInput),
    .io_addInput(mac_20_6_io_addInput),
    .io_output(mac_20_6_io_output),
    .io_passthrough(mac_20_6_io_passthrough)
  );
  MAC mac_20_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_7_clock),
    .reset(mac_20_7_reset),
    .io_load(mac_20_7_io_load),
    .io_mulInput(mac_20_7_io_mulInput),
    .io_addInput(mac_20_7_io_addInput),
    .io_output(mac_20_7_io_output),
    .io_passthrough(mac_20_7_io_passthrough)
  );
  MAC mac_20_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_8_clock),
    .reset(mac_20_8_reset),
    .io_load(mac_20_8_io_load),
    .io_mulInput(mac_20_8_io_mulInput),
    .io_addInput(mac_20_8_io_addInput),
    .io_output(mac_20_8_io_output),
    .io_passthrough(mac_20_8_io_passthrough)
  );
  MAC mac_20_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_9_clock),
    .reset(mac_20_9_reset),
    .io_load(mac_20_9_io_load),
    .io_mulInput(mac_20_9_io_mulInput),
    .io_addInput(mac_20_9_io_addInput),
    .io_output(mac_20_9_io_output),
    .io_passthrough(mac_20_9_io_passthrough)
  );
  MAC mac_20_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_10_clock),
    .reset(mac_20_10_reset),
    .io_load(mac_20_10_io_load),
    .io_mulInput(mac_20_10_io_mulInput),
    .io_addInput(mac_20_10_io_addInput),
    .io_output(mac_20_10_io_output),
    .io_passthrough(mac_20_10_io_passthrough)
  );
  MAC mac_20_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_11_clock),
    .reset(mac_20_11_reset),
    .io_load(mac_20_11_io_load),
    .io_mulInput(mac_20_11_io_mulInput),
    .io_addInput(mac_20_11_io_addInput),
    .io_output(mac_20_11_io_output),
    .io_passthrough(mac_20_11_io_passthrough)
  );
  MAC mac_20_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_12_clock),
    .reset(mac_20_12_reset),
    .io_load(mac_20_12_io_load),
    .io_mulInput(mac_20_12_io_mulInput),
    .io_addInput(mac_20_12_io_addInput),
    .io_output(mac_20_12_io_output),
    .io_passthrough(mac_20_12_io_passthrough)
  );
  MAC mac_20_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_13_clock),
    .reset(mac_20_13_reset),
    .io_load(mac_20_13_io_load),
    .io_mulInput(mac_20_13_io_mulInput),
    .io_addInput(mac_20_13_io_addInput),
    .io_output(mac_20_13_io_output),
    .io_passthrough(mac_20_13_io_passthrough)
  );
  MAC mac_20_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_14_clock),
    .reset(mac_20_14_reset),
    .io_load(mac_20_14_io_load),
    .io_mulInput(mac_20_14_io_mulInput),
    .io_addInput(mac_20_14_io_addInput),
    .io_output(mac_20_14_io_output),
    .io_passthrough(mac_20_14_io_passthrough)
  );
  MAC mac_20_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_15_clock),
    .reset(mac_20_15_reset),
    .io_load(mac_20_15_io_load),
    .io_mulInput(mac_20_15_io_mulInput),
    .io_addInput(mac_20_15_io_addInput),
    .io_output(mac_20_15_io_output),
    .io_passthrough(mac_20_15_io_passthrough)
  );
  MAC mac_20_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_16_clock),
    .reset(mac_20_16_reset),
    .io_load(mac_20_16_io_load),
    .io_mulInput(mac_20_16_io_mulInput),
    .io_addInput(mac_20_16_io_addInput),
    .io_output(mac_20_16_io_output),
    .io_passthrough(mac_20_16_io_passthrough)
  );
  MAC mac_20_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_17_clock),
    .reset(mac_20_17_reset),
    .io_load(mac_20_17_io_load),
    .io_mulInput(mac_20_17_io_mulInput),
    .io_addInput(mac_20_17_io_addInput),
    .io_output(mac_20_17_io_output),
    .io_passthrough(mac_20_17_io_passthrough)
  );
  MAC mac_20_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_18_clock),
    .reset(mac_20_18_reset),
    .io_load(mac_20_18_io_load),
    .io_mulInput(mac_20_18_io_mulInput),
    .io_addInput(mac_20_18_io_addInput),
    .io_output(mac_20_18_io_output),
    .io_passthrough(mac_20_18_io_passthrough)
  );
  MAC mac_20_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_19_clock),
    .reset(mac_20_19_reset),
    .io_load(mac_20_19_io_load),
    .io_mulInput(mac_20_19_io_mulInput),
    .io_addInput(mac_20_19_io_addInput),
    .io_output(mac_20_19_io_output),
    .io_passthrough(mac_20_19_io_passthrough)
  );
  MAC mac_20_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_20_clock),
    .reset(mac_20_20_reset),
    .io_load(mac_20_20_io_load),
    .io_mulInput(mac_20_20_io_mulInput),
    .io_addInput(mac_20_20_io_addInput),
    .io_output(mac_20_20_io_output),
    .io_passthrough(mac_20_20_io_passthrough)
  );
  MAC mac_20_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_21_clock),
    .reset(mac_20_21_reset),
    .io_load(mac_20_21_io_load),
    .io_mulInput(mac_20_21_io_mulInput),
    .io_addInput(mac_20_21_io_addInput),
    .io_output(mac_20_21_io_output),
    .io_passthrough(mac_20_21_io_passthrough)
  );
  MAC mac_20_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_22_clock),
    .reset(mac_20_22_reset),
    .io_load(mac_20_22_io_load),
    .io_mulInput(mac_20_22_io_mulInput),
    .io_addInput(mac_20_22_io_addInput),
    .io_output(mac_20_22_io_output),
    .io_passthrough(mac_20_22_io_passthrough)
  );
  MAC mac_20_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_23_clock),
    .reset(mac_20_23_reset),
    .io_load(mac_20_23_io_load),
    .io_mulInput(mac_20_23_io_mulInput),
    .io_addInput(mac_20_23_io_addInput),
    .io_output(mac_20_23_io_output),
    .io_passthrough(mac_20_23_io_passthrough)
  );
  MAC mac_20_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_24_clock),
    .reset(mac_20_24_reset),
    .io_load(mac_20_24_io_load),
    .io_mulInput(mac_20_24_io_mulInput),
    .io_addInput(mac_20_24_io_addInput),
    .io_output(mac_20_24_io_output),
    .io_passthrough(mac_20_24_io_passthrough)
  );
  MAC mac_20_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_25_clock),
    .reset(mac_20_25_reset),
    .io_load(mac_20_25_io_load),
    .io_mulInput(mac_20_25_io_mulInput),
    .io_addInput(mac_20_25_io_addInput),
    .io_output(mac_20_25_io_output),
    .io_passthrough(mac_20_25_io_passthrough)
  );
  MAC mac_20_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_26_clock),
    .reset(mac_20_26_reset),
    .io_load(mac_20_26_io_load),
    .io_mulInput(mac_20_26_io_mulInput),
    .io_addInput(mac_20_26_io_addInput),
    .io_output(mac_20_26_io_output),
    .io_passthrough(mac_20_26_io_passthrough)
  );
  MAC mac_20_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_27_clock),
    .reset(mac_20_27_reset),
    .io_load(mac_20_27_io_load),
    .io_mulInput(mac_20_27_io_mulInput),
    .io_addInput(mac_20_27_io_addInput),
    .io_output(mac_20_27_io_output),
    .io_passthrough(mac_20_27_io_passthrough)
  );
  MAC mac_20_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_28_clock),
    .reset(mac_20_28_reset),
    .io_load(mac_20_28_io_load),
    .io_mulInput(mac_20_28_io_mulInput),
    .io_addInput(mac_20_28_io_addInput),
    .io_output(mac_20_28_io_output),
    .io_passthrough(mac_20_28_io_passthrough)
  );
  MAC mac_20_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_29_clock),
    .reset(mac_20_29_reset),
    .io_load(mac_20_29_io_load),
    .io_mulInput(mac_20_29_io_mulInput),
    .io_addInput(mac_20_29_io_addInput),
    .io_output(mac_20_29_io_output),
    .io_passthrough(mac_20_29_io_passthrough)
  );
  MAC mac_20_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_30_clock),
    .reset(mac_20_30_reset),
    .io_load(mac_20_30_io_load),
    .io_mulInput(mac_20_30_io_mulInput),
    .io_addInput(mac_20_30_io_addInput),
    .io_output(mac_20_30_io_output),
    .io_passthrough(mac_20_30_io_passthrough)
  );
  MAC mac_20_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_20_31_clock),
    .reset(mac_20_31_reset),
    .io_load(mac_20_31_io_load),
    .io_mulInput(mac_20_31_io_mulInput),
    .io_addInput(mac_20_31_io_addInput),
    .io_output(mac_20_31_io_output),
    .io_passthrough(mac_20_31_io_passthrough)
  );
  MAC mac_21_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_0_clock),
    .reset(mac_21_0_reset),
    .io_load(mac_21_0_io_load),
    .io_mulInput(mac_21_0_io_mulInput),
    .io_addInput(mac_21_0_io_addInput),
    .io_output(mac_21_0_io_output),
    .io_passthrough(mac_21_0_io_passthrough)
  );
  MAC mac_21_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_1_clock),
    .reset(mac_21_1_reset),
    .io_load(mac_21_1_io_load),
    .io_mulInput(mac_21_1_io_mulInput),
    .io_addInput(mac_21_1_io_addInput),
    .io_output(mac_21_1_io_output),
    .io_passthrough(mac_21_1_io_passthrough)
  );
  MAC mac_21_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_2_clock),
    .reset(mac_21_2_reset),
    .io_load(mac_21_2_io_load),
    .io_mulInput(mac_21_2_io_mulInput),
    .io_addInput(mac_21_2_io_addInput),
    .io_output(mac_21_2_io_output),
    .io_passthrough(mac_21_2_io_passthrough)
  );
  MAC mac_21_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_3_clock),
    .reset(mac_21_3_reset),
    .io_load(mac_21_3_io_load),
    .io_mulInput(mac_21_3_io_mulInput),
    .io_addInput(mac_21_3_io_addInput),
    .io_output(mac_21_3_io_output),
    .io_passthrough(mac_21_3_io_passthrough)
  );
  MAC mac_21_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_4_clock),
    .reset(mac_21_4_reset),
    .io_load(mac_21_4_io_load),
    .io_mulInput(mac_21_4_io_mulInput),
    .io_addInput(mac_21_4_io_addInput),
    .io_output(mac_21_4_io_output),
    .io_passthrough(mac_21_4_io_passthrough)
  );
  MAC mac_21_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_5_clock),
    .reset(mac_21_5_reset),
    .io_load(mac_21_5_io_load),
    .io_mulInput(mac_21_5_io_mulInput),
    .io_addInput(mac_21_5_io_addInput),
    .io_output(mac_21_5_io_output),
    .io_passthrough(mac_21_5_io_passthrough)
  );
  MAC mac_21_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_6_clock),
    .reset(mac_21_6_reset),
    .io_load(mac_21_6_io_load),
    .io_mulInput(mac_21_6_io_mulInput),
    .io_addInput(mac_21_6_io_addInput),
    .io_output(mac_21_6_io_output),
    .io_passthrough(mac_21_6_io_passthrough)
  );
  MAC mac_21_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_7_clock),
    .reset(mac_21_7_reset),
    .io_load(mac_21_7_io_load),
    .io_mulInput(mac_21_7_io_mulInput),
    .io_addInput(mac_21_7_io_addInput),
    .io_output(mac_21_7_io_output),
    .io_passthrough(mac_21_7_io_passthrough)
  );
  MAC mac_21_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_8_clock),
    .reset(mac_21_8_reset),
    .io_load(mac_21_8_io_load),
    .io_mulInput(mac_21_8_io_mulInput),
    .io_addInput(mac_21_8_io_addInput),
    .io_output(mac_21_8_io_output),
    .io_passthrough(mac_21_8_io_passthrough)
  );
  MAC mac_21_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_9_clock),
    .reset(mac_21_9_reset),
    .io_load(mac_21_9_io_load),
    .io_mulInput(mac_21_9_io_mulInput),
    .io_addInput(mac_21_9_io_addInput),
    .io_output(mac_21_9_io_output),
    .io_passthrough(mac_21_9_io_passthrough)
  );
  MAC mac_21_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_10_clock),
    .reset(mac_21_10_reset),
    .io_load(mac_21_10_io_load),
    .io_mulInput(mac_21_10_io_mulInput),
    .io_addInput(mac_21_10_io_addInput),
    .io_output(mac_21_10_io_output),
    .io_passthrough(mac_21_10_io_passthrough)
  );
  MAC mac_21_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_11_clock),
    .reset(mac_21_11_reset),
    .io_load(mac_21_11_io_load),
    .io_mulInput(mac_21_11_io_mulInput),
    .io_addInput(mac_21_11_io_addInput),
    .io_output(mac_21_11_io_output),
    .io_passthrough(mac_21_11_io_passthrough)
  );
  MAC mac_21_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_12_clock),
    .reset(mac_21_12_reset),
    .io_load(mac_21_12_io_load),
    .io_mulInput(mac_21_12_io_mulInput),
    .io_addInput(mac_21_12_io_addInput),
    .io_output(mac_21_12_io_output),
    .io_passthrough(mac_21_12_io_passthrough)
  );
  MAC mac_21_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_13_clock),
    .reset(mac_21_13_reset),
    .io_load(mac_21_13_io_load),
    .io_mulInput(mac_21_13_io_mulInput),
    .io_addInput(mac_21_13_io_addInput),
    .io_output(mac_21_13_io_output),
    .io_passthrough(mac_21_13_io_passthrough)
  );
  MAC mac_21_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_14_clock),
    .reset(mac_21_14_reset),
    .io_load(mac_21_14_io_load),
    .io_mulInput(mac_21_14_io_mulInput),
    .io_addInput(mac_21_14_io_addInput),
    .io_output(mac_21_14_io_output),
    .io_passthrough(mac_21_14_io_passthrough)
  );
  MAC mac_21_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_15_clock),
    .reset(mac_21_15_reset),
    .io_load(mac_21_15_io_load),
    .io_mulInput(mac_21_15_io_mulInput),
    .io_addInput(mac_21_15_io_addInput),
    .io_output(mac_21_15_io_output),
    .io_passthrough(mac_21_15_io_passthrough)
  );
  MAC mac_21_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_16_clock),
    .reset(mac_21_16_reset),
    .io_load(mac_21_16_io_load),
    .io_mulInput(mac_21_16_io_mulInput),
    .io_addInput(mac_21_16_io_addInput),
    .io_output(mac_21_16_io_output),
    .io_passthrough(mac_21_16_io_passthrough)
  );
  MAC mac_21_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_17_clock),
    .reset(mac_21_17_reset),
    .io_load(mac_21_17_io_load),
    .io_mulInput(mac_21_17_io_mulInput),
    .io_addInput(mac_21_17_io_addInput),
    .io_output(mac_21_17_io_output),
    .io_passthrough(mac_21_17_io_passthrough)
  );
  MAC mac_21_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_18_clock),
    .reset(mac_21_18_reset),
    .io_load(mac_21_18_io_load),
    .io_mulInput(mac_21_18_io_mulInput),
    .io_addInput(mac_21_18_io_addInput),
    .io_output(mac_21_18_io_output),
    .io_passthrough(mac_21_18_io_passthrough)
  );
  MAC mac_21_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_19_clock),
    .reset(mac_21_19_reset),
    .io_load(mac_21_19_io_load),
    .io_mulInput(mac_21_19_io_mulInput),
    .io_addInput(mac_21_19_io_addInput),
    .io_output(mac_21_19_io_output),
    .io_passthrough(mac_21_19_io_passthrough)
  );
  MAC mac_21_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_20_clock),
    .reset(mac_21_20_reset),
    .io_load(mac_21_20_io_load),
    .io_mulInput(mac_21_20_io_mulInput),
    .io_addInput(mac_21_20_io_addInput),
    .io_output(mac_21_20_io_output),
    .io_passthrough(mac_21_20_io_passthrough)
  );
  MAC mac_21_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_21_clock),
    .reset(mac_21_21_reset),
    .io_load(mac_21_21_io_load),
    .io_mulInput(mac_21_21_io_mulInput),
    .io_addInput(mac_21_21_io_addInput),
    .io_output(mac_21_21_io_output),
    .io_passthrough(mac_21_21_io_passthrough)
  );
  MAC mac_21_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_22_clock),
    .reset(mac_21_22_reset),
    .io_load(mac_21_22_io_load),
    .io_mulInput(mac_21_22_io_mulInput),
    .io_addInput(mac_21_22_io_addInput),
    .io_output(mac_21_22_io_output),
    .io_passthrough(mac_21_22_io_passthrough)
  );
  MAC mac_21_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_23_clock),
    .reset(mac_21_23_reset),
    .io_load(mac_21_23_io_load),
    .io_mulInput(mac_21_23_io_mulInput),
    .io_addInput(mac_21_23_io_addInput),
    .io_output(mac_21_23_io_output),
    .io_passthrough(mac_21_23_io_passthrough)
  );
  MAC mac_21_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_24_clock),
    .reset(mac_21_24_reset),
    .io_load(mac_21_24_io_load),
    .io_mulInput(mac_21_24_io_mulInput),
    .io_addInput(mac_21_24_io_addInput),
    .io_output(mac_21_24_io_output),
    .io_passthrough(mac_21_24_io_passthrough)
  );
  MAC mac_21_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_25_clock),
    .reset(mac_21_25_reset),
    .io_load(mac_21_25_io_load),
    .io_mulInput(mac_21_25_io_mulInput),
    .io_addInput(mac_21_25_io_addInput),
    .io_output(mac_21_25_io_output),
    .io_passthrough(mac_21_25_io_passthrough)
  );
  MAC mac_21_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_26_clock),
    .reset(mac_21_26_reset),
    .io_load(mac_21_26_io_load),
    .io_mulInput(mac_21_26_io_mulInput),
    .io_addInput(mac_21_26_io_addInput),
    .io_output(mac_21_26_io_output),
    .io_passthrough(mac_21_26_io_passthrough)
  );
  MAC mac_21_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_27_clock),
    .reset(mac_21_27_reset),
    .io_load(mac_21_27_io_load),
    .io_mulInput(mac_21_27_io_mulInput),
    .io_addInput(mac_21_27_io_addInput),
    .io_output(mac_21_27_io_output),
    .io_passthrough(mac_21_27_io_passthrough)
  );
  MAC mac_21_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_28_clock),
    .reset(mac_21_28_reset),
    .io_load(mac_21_28_io_load),
    .io_mulInput(mac_21_28_io_mulInput),
    .io_addInput(mac_21_28_io_addInput),
    .io_output(mac_21_28_io_output),
    .io_passthrough(mac_21_28_io_passthrough)
  );
  MAC mac_21_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_29_clock),
    .reset(mac_21_29_reset),
    .io_load(mac_21_29_io_load),
    .io_mulInput(mac_21_29_io_mulInput),
    .io_addInput(mac_21_29_io_addInput),
    .io_output(mac_21_29_io_output),
    .io_passthrough(mac_21_29_io_passthrough)
  );
  MAC mac_21_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_30_clock),
    .reset(mac_21_30_reset),
    .io_load(mac_21_30_io_load),
    .io_mulInput(mac_21_30_io_mulInput),
    .io_addInput(mac_21_30_io_addInput),
    .io_output(mac_21_30_io_output),
    .io_passthrough(mac_21_30_io_passthrough)
  );
  MAC mac_21_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_21_31_clock),
    .reset(mac_21_31_reset),
    .io_load(mac_21_31_io_load),
    .io_mulInput(mac_21_31_io_mulInput),
    .io_addInput(mac_21_31_io_addInput),
    .io_output(mac_21_31_io_output),
    .io_passthrough(mac_21_31_io_passthrough)
  );
  MAC mac_22_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_0_clock),
    .reset(mac_22_0_reset),
    .io_load(mac_22_0_io_load),
    .io_mulInput(mac_22_0_io_mulInput),
    .io_addInput(mac_22_0_io_addInput),
    .io_output(mac_22_0_io_output),
    .io_passthrough(mac_22_0_io_passthrough)
  );
  MAC mac_22_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_1_clock),
    .reset(mac_22_1_reset),
    .io_load(mac_22_1_io_load),
    .io_mulInput(mac_22_1_io_mulInput),
    .io_addInput(mac_22_1_io_addInput),
    .io_output(mac_22_1_io_output),
    .io_passthrough(mac_22_1_io_passthrough)
  );
  MAC mac_22_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_2_clock),
    .reset(mac_22_2_reset),
    .io_load(mac_22_2_io_load),
    .io_mulInput(mac_22_2_io_mulInput),
    .io_addInput(mac_22_2_io_addInput),
    .io_output(mac_22_2_io_output),
    .io_passthrough(mac_22_2_io_passthrough)
  );
  MAC mac_22_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_3_clock),
    .reset(mac_22_3_reset),
    .io_load(mac_22_3_io_load),
    .io_mulInput(mac_22_3_io_mulInput),
    .io_addInput(mac_22_3_io_addInput),
    .io_output(mac_22_3_io_output),
    .io_passthrough(mac_22_3_io_passthrough)
  );
  MAC mac_22_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_4_clock),
    .reset(mac_22_4_reset),
    .io_load(mac_22_4_io_load),
    .io_mulInput(mac_22_4_io_mulInput),
    .io_addInput(mac_22_4_io_addInput),
    .io_output(mac_22_4_io_output),
    .io_passthrough(mac_22_4_io_passthrough)
  );
  MAC mac_22_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_5_clock),
    .reset(mac_22_5_reset),
    .io_load(mac_22_5_io_load),
    .io_mulInput(mac_22_5_io_mulInput),
    .io_addInput(mac_22_5_io_addInput),
    .io_output(mac_22_5_io_output),
    .io_passthrough(mac_22_5_io_passthrough)
  );
  MAC mac_22_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_6_clock),
    .reset(mac_22_6_reset),
    .io_load(mac_22_6_io_load),
    .io_mulInput(mac_22_6_io_mulInput),
    .io_addInput(mac_22_6_io_addInput),
    .io_output(mac_22_6_io_output),
    .io_passthrough(mac_22_6_io_passthrough)
  );
  MAC mac_22_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_7_clock),
    .reset(mac_22_7_reset),
    .io_load(mac_22_7_io_load),
    .io_mulInput(mac_22_7_io_mulInput),
    .io_addInput(mac_22_7_io_addInput),
    .io_output(mac_22_7_io_output),
    .io_passthrough(mac_22_7_io_passthrough)
  );
  MAC mac_22_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_8_clock),
    .reset(mac_22_8_reset),
    .io_load(mac_22_8_io_load),
    .io_mulInput(mac_22_8_io_mulInput),
    .io_addInput(mac_22_8_io_addInput),
    .io_output(mac_22_8_io_output),
    .io_passthrough(mac_22_8_io_passthrough)
  );
  MAC mac_22_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_9_clock),
    .reset(mac_22_9_reset),
    .io_load(mac_22_9_io_load),
    .io_mulInput(mac_22_9_io_mulInput),
    .io_addInput(mac_22_9_io_addInput),
    .io_output(mac_22_9_io_output),
    .io_passthrough(mac_22_9_io_passthrough)
  );
  MAC mac_22_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_10_clock),
    .reset(mac_22_10_reset),
    .io_load(mac_22_10_io_load),
    .io_mulInput(mac_22_10_io_mulInput),
    .io_addInput(mac_22_10_io_addInput),
    .io_output(mac_22_10_io_output),
    .io_passthrough(mac_22_10_io_passthrough)
  );
  MAC mac_22_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_11_clock),
    .reset(mac_22_11_reset),
    .io_load(mac_22_11_io_load),
    .io_mulInput(mac_22_11_io_mulInput),
    .io_addInput(mac_22_11_io_addInput),
    .io_output(mac_22_11_io_output),
    .io_passthrough(mac_22_11_io_passthrough)
  );
  MAC mac_22_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_12_clock),
    .reset(mac_22_12_reset),
    .io_load(mac_22_12_io_load),
    .io_mulInput(mac_22_12_io_mulInput),
    .io_addInput(mac_22_12_io_addInput),
    .io_output(mac_22_12_io_output),
    .io_passthrough(mac_22_12_io_passthrough)
  );
  MAC mac_22_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_13_clock),
    .reset(mac_22_13_reset),
    .io_load(mac_22_13_io_load),
    .io_mulInput(mac_22_13_io_mulInput),
    .io_addInput(mac_22_13_io_addInput),
    .io_output(mac_22_13_io_output),
    .io_passthrough(mac_22_13_io_passthrough)
  );
  MAC mac_22_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_14_clock),
    .reset(mac_22_14_reset),
    .io_load(mac_22_14_io_load),
    .io_mulInput(mac_22_14_io_mulInput),
    .io_addInput(mac_22_14_io_addInput),
    .io_output(mac_22_14_io_output),
    .io_passthrough(mac_22_14_io_passthrough)
  );
  MAC mac_22_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_15_clock),
    .reset(mac_22_15_reset),
    .io_load(mac_22_15_io_load),
    .io_mulInput(mac_22_15_io_mulInput),
    .io_addInput(mac_22_15_io_addInput),
    .io_output(mac_22_15_io_output),
    .io_passthrough(mac_22_15_io_passthrough)
  );
  MAC mac_22_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_16_clock),
    .reset(mac_22_16_reset),
    .io_load(mac_22_16_io_load),
    .io_mulInput(mac_22_16_io_mulInput),
    .io_addInput(mac_22_16_io_addInput),
    .io_output(mac_22_16_io_output),
    .io_passthrough(mac_22_16_io_passthrough)
  );
  MAC mac_22_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_17_clock),
    .reset(mac_22_17_reset),
    .io_load(mac_22_17_io_load),
    .io_mulInput(mac_22_17_io_mulInput),
    .io_addInput(mac_22_17_io_addInput),
    .io_output(mac_22_17_io_output),
    .io_passthrough(mac_22_17_io_passthrough)
  );
  MAC mac_22_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_18_clock),
    .reset(mac_22_18_reset),
    .io_load(mac_22_18_io_load),
    .io_mulInput(mac_22_18_io_mulInput),
    .io_addInput(mac_22_18_io_addInput),
    .io_output(mac_22_18_io_output),
    .io_passthrough(mac_22_18_io_passthrough)
  );
  MAC mac_22_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_19_clock),
    .reset(mac_22_19_reset),
    .io_load(mac_22_19_io_load),
    .io_mulInput(mac_22_19_io_mulInput),
    .io_addInput(mac_22_19_io_addInput),
    .io_output(mac_22_19_io_output),
    .io_passthrough(mac_22_19_io_passthrough)
  );
  MAC mac_22_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_20_clock),
    .reset(mac_22_20_reset),
    .io_load(mac_22_20_io_load),
    .io_mulInput(mac_22_20_io_mulInput),
    .io_addInput(mac_22_20_io_addInput),
    .io_output(mac_22_20_io_output),
    .io_passthrough(mac_22_20_io_passthrough)
  );
  MAC mac_22_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_21_clock),
    .reset(mac_22_21_reset),
    .io_load(mac_22_21_io_load),
    .io_mulInput(mac_22_21_io_mulInput),
    .io_addInput(mac_22_21_io_addInput),
    .io_output(mac_22_21_io_output),
    .io_passthrough(mac_22_21_io_passthrough)
  );
  MAC mac_22_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_22_clock),
    .reset(mac_22_22_reset),
    .io_load(mac_22_22_io_load),
    .io_mulInput(mac_22_22_io_mulInput),
    .io_addInput(mac_22_22_io_addInput),
    .io_output(mac_22_22_io_output),
    .io_passthrough(mac_22_22_io_passthrough)
  );
  MAC mac_22_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_23_clock),
    .reset(mac_22_23_reset),
    .io_load(mac_22_23_io_load),
    .io_mulInput(mac_22_23_io_mulInput),
    .io_addInput(mac_22_23_io_addInput),
    .io_output(mac_22_23_io_output),
    .io_passthrough(mac_22_23_io_passthrough)
  );
  MAC mac_22_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_24_clock),
    .reset(mac_22_24_reset),
    .io_load(mac_22_24_io_load),
    .io_mulInput(mac_22_24_io_mulInput),
    .io_addInput(mac_22_24_io_addInput),
    .io_output(mac_22_24_io_output),
    .io_passthrough(mac_22_24_io_passthrough)
  );
  MAC mac_22_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_25_clock),
    .reset(mac_22_25_reset),
    .io_load(mac_22_25_io_load),
    .io_mulInput(mac_22_25_io_mulInput),
    .io_addInput(mac_22_25_io_addInput),
    .io_output(mac_22_25_io_output),
    .io_passthrough(mac_22_25_io_passthrough)
  );
  MAC mac_22_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_26_clock),
    .reset(mac_22_26_reset),
    .io_load(mac_22_26_io_load),
    .io_mulInput(mac_22_26_io_mulInput),
    .io_addInput(mac_22_26_io_addInput),
    .io_output(mac_22_26_io_output),
    .io_passthrough(mac_22_26_io_passthrough)
  );
  MAC mac_22_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_27_clock),
    .reset(mac_22_27_reset),
    .io_load(mac_22_27_io_load),
    .io_mulInput(mac_22_27_io_mulInput),
    .io_addInput(mac_22_27_io_addInput),
    .io_output(mac_22_27_io_output),
    .io_passthrough(mac_22_27_io_passthrough)
  );
  MAC mac_22_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_28_clock),
    .reset(mac_22_28_reset),
    .io_load(mac_22_28_io_load),
    .io_mulInput(mac_22_28_io_mulInput),
    .io_addInput(mac_22_28_io_addInput),
    .io_output(mac_22_28_io_output),
    .io_passthrough(mac_22_28_io_passthrough)
  );
  MAC mac_22_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_29_clock),
    .reset(mac_22_29_reset),
    .io_load(mac_22_29_io_load),
    .io_mulInput(mac_22_29_io_mulInput),
    .io_addInput(mac_22_29_io_addInput),
    .io_output(mac_22_29_io_output),
    .io_passthrough(mac_22_29_io_passthrough)
  );
  MAC mac_22_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_30_clock),
    .reset(mac_22_30_reset),
    .io_load(mac_22_30_io_load),
    .io_mulInput(mac_22_30_io_mulInput),
    .io_addInput(mac_22_30_io_addInput),
    .io_output(mac_22_30_io_output),
    .io_passthrough(mac_22_30_io_passthrough)
  );
  MAC mac_22_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_22_31_clock),
    .reset(mac_22_31_reset),
    .io_load(mac_22_31_io_load),
    .io_mulInput(mac_22_31_io_mulInput),
    .io_addInput(mac_22_31_io_addInput),
    .io_output(mac_22_31_io_output),
    .io_passthrough(mac_22_31_io_passthrough)
  );
  MAC mac_23_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_0_clock),
    .reset(mac_23_0_reset),
    .io_load(mac_23_0_io_load),
    .io_mulInput(mac_23_0_io_mulInput),
    .io_addInput(mac_23_0_io_addInput),
    .io_output(mac_23_0_io_output),
    .io_passthrough(mac_23_0_io_passthrough)
  );
  MAC mac_23_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_1_clock),
    .reset(mac_23_1_reset),
    .io_load(mac_23_1_io_load),
    .io_mulInput(mac_23_1_io_mulInput),
    .io_addInput(mac_23_1_io_addInput),
    .io_output(mac_23_1_io_output),
    .io_passthrough(mac_23_1_io_passthrough)
  );
  MAC mac_23_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_2_clock),
    .reset(mac_23_2_reset),
    .io_load(mac_23_2_io_load),
    .io_mulInput(mac_23_2_io_mulInput),
    .io_addInput(mac_23_2_io_addInput),
    .io_output(mac_23_2_io_output),
    .io_passthrough(mac_23_2_io_passthrough)
  );
  MAC mac_23_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_3_clock),
    .reset(mac_23_3_reset),
    .io_load(mac_23_3_io_load),
    .io_mulInput(mac_23_3_io_mulInput),
    .io_addInput(mac_23_3_io_addInput),
    .io_output(mac_23_3_io_output),
    .io_passthrough(mac_23_3_io_passthrough)
  );
  MAC mac_23_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_4_clock),
    .reset(mac_23_4_reset),
    .io_load(mac_23_4_io_load),
    .io_mulInput(mac_23_4_io_mulInput),
    .io_addInput(mac_23_4_io_addInput),
    .io_output(mac_23_4_io_output),
    .io_passthrough(mac_23_4_io_passthrough)
  );
  MAC mac_23_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_5_clock),
    .reset(mac_23_5_reset),
    .io_load(mac_23_5_io_load),
    .io_mulInput(mac_23_5_io_mulInput),
    .io_addInput(mac_23_5_io_addInput),
    .io_output(mac_23_5_io_output),
    .io_passthrough(mac_23_5_io_passthrough)
  );
  MAC mac_23_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_6_clock),
    .reset(mac_23_6_reset),
    .io_load(mac_23_6_io_load),
    .io_mulInput(mac_23_6_io_mulInput),
    .io_addInput(mac_23_6_io_addInput),
    .io_output(mac_23_6_io_output),
    .io_passthrough(mac_23_6_io_passthrough)
  );
  MAC mac_23_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_7_clock),
    .reset(mac_23_7_reset),
    .io_load(mac_23_7_io_load),
    .io_mulInput(mac_23_7_io_mulInput),
    .io_addInput(mac_23_7_io_addInput),
    .io_output(mac_23_7_io_output),
    .io_passthrough(mac_23_7_io_passthrough)
  );
  MAC mac_23_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_8_clock),
    .reset(mac_23_8_reset),
    .io_load(mac_23_8_io_load),
    .io_mulInput(mac_23_8_io_mulInput),
    .io_addInput(mac_23_8_io_addInput),
    .io_output(mac_23_8_io_output),
    .io_passthrough(mac_23_8_io_passthrough)
  );
  MAC mac_23_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_9_clock),
    .reset(mac_23_9_reset),
    .io_load(mac_23_9_io_load),
    .io_mulInput(mac_23_9_io_mulInput),
    .io_addInput(mac_23_9_io_addInput),
    .io_output(mac_23_9_io_output),
    .io_passthrough(mac_23_9_io_passthrough)
  );
  MAC mac_23_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_10_clock),
    .reset(mac_23_10_reset),
    .io_load(mac_23_10_io_load),
    .io_mulInput(mac_23_10_io_mulInput),
    .io_addInput(mac_23_10_io_addInput),
    .io_output(mac_23_10_io_output),
    .io_passthrough(mac_23_10_io_passthrough)
  );
  MAC mac_23_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_11_clock),
    .reset(mac_23_11_reset),
    .io_load(mac_23_11_io_load),
    .io_mulInput(mac_23_11_io_mulInput),
    .io_addInput(mac_23_11_io_addInput),
    .io_output(mac_23_11_io_output),
    .io_passthrough(mac_23_11_io_passthrough)
  );
  MAC mac_23_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_12_clock),
    .reset(mac_23_12_reset),
    .io_load(mac_23_12_io_load),
    .io_mulInput(mac_23_12_io_mulInput),
    .io_addInput(mac_23_12_io_addInput),
    .io_output(mac_23_12_io_output),
    .io_passthrough(mac_23_12_io_passthrough)
  );
  MAC mac_23_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_13_clock),
    .reset(mac_23_13_reset),
    .io_load(mac_23_13_io_load),
    .io_mulInput(mac_23_13_io_mulInput),
    .io_addInput(mac_23_13_io_addInput),
    .io_output(mac_23_13_io_output),
    .io_passthrough(mac_23_13_io_passthrough)
  );
  MAC mac_23_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_14_clock),
    .reset(mac_23_14_reset),
    .io_load(mac_23_14_io_load),
    .io_mulInput(mac_23_14_io_mulInput),
    .io_addInput(mac_23_14_io_addInput),
    .io_output(mac_23_14_io_output),
    .io_passthrough(mac_23_14_io_passthrough)
  );
  MAC mac_23_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_15_clock),
    .reset(mac_23_15_reset),
    .io_load(mac_23_15_io_load),
    .io_mulInput(mac_23_15_io_mulInput),
    .io_addInput(mac_23_15_io_addInput),
    .io_output(mac_23_15_io_output),
    .io_passthrough(mac_23_15_io_passthrough)
  );
  MAC mac_23_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_16_clock),
    .reset(mac_23_16_reset),
    .io_load(mac_23_16_io_load),
    .io_mulInput(mac_23_16_io_mulInput),
    .io_addInput(mac_23_16_io_addInput),
    .io_output(mac_23_16_io_output),
    .io_passthrough(mac_23_16_io_passthrough)
  );
  MAC mac_23_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_17_clock),
    .reset(mac_23_17_reset),
    .io_load(mac_23_17_io_load),
    .io_mulInput(mac_23_17_io_mulInput),
    .io_addInput(mac_23_17_io_addInput),
    .io_output(mac_23_17_io_output),
    .io_passthrough(mac_23_17_io_passthrough)
  );
  MAC mac_23_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_18_clock),
    .reset(mac_23_18_reset),
    .io_load(mac_23_18_io_load),
    .io_mulInput(mac_23_18_io_mulInput),
    .io_addInput(mac_23_18_io_addInput),
    .io_output(mac_23_18_io_output),
    .io_passthrough(mac_23_18_io_passthrough)
  );
  MAC mac_23_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_19_clock),
    .reset(mac_23_19_reset),
    .io_load(mac_23_19_io_load),
    .io_mulInput(mac_23_19_io_mulInput),
    .io_addInput(mac_23_19_io_addInput),
    .io_output(mac_23_19_io_output),
    .io_passthrough(mac_23_19_io_passthrough)
  );
  MAC mac_23_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_20_clock),
    .reset(mac_23_20_reset),
    .io_load(mac_23_20_io_load),
    .io_mulInput(mac_23_20_io_mulInput),
    .io_addInput(mac_23_20_io_addInput),
    .io_output(mac_23_20_io_output),
    .io_passthrough(mac_23_20_io_passthrough)
  );
  MAC mac_23_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_21_clock),
    .reset(mac_23_21_reset),
    .io_load(mac_23_21_io_load),
    .io_mulInput(mac_23_21_io_mulInput),
    .io_addInput(mac_23_21_io_addInput),
    .io_output(mac_23_21_io_output),
    .io_passthrough(mac_23_21_io_passthrough)
  );
  MAC mac_23_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_22_clock),
    .reset(mac_23_22_reset),
    .io_load(mac_23_22_io_load),
    .io_mulInput(mac_23_22_io_mulInput),
    .io_addInput(mac_23_22_io_addInput),
    .io_output(mac_23_22_io_output),
    .io_passthrough(mac_23_22_io_passthrough)
  );
  MAC mac_23_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_23_clock),
    .reset(mac_23_23_reset),
    .io_load(mac_23_23_io_load),
    .io_mulInput(mac_23_23_io_mulInput),
    .io_addInput(mac_23_23_io_addInput),
    .io_output(mac_23_23_io_output),
    .io_passthrough(mac_23_23_io_passthrough)
  );
  MAC mac_23_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_24_clock),
    .reset(mac_23_24_reset),
    .io_load(mac_23_24_io_load),
    .io_mulInput(mac_23_24_io_mulInput),
    .io_addInput(mac_23_24_io_addInput),
    .io_output(mac_23_24_io_output),
    .io_passthrough(mac_23_24_io_passthrough)
  );
  MAC mac_23_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_25_clock),
    .reset(mac_23_25_reset),
    .io_load(mac_23_25_io_load),
    .io_mulInput(mac_23_25_io_mulInput),
    .io_addInput(mac_23_25_io_addInput),
    .io_output(mac_23_25_io_output),
    .io_passthrough(mac_23_25_io_passthrough)
  );
  MAC mac_23_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_26_clock),
    .reset(mac_23_26_reset),
    .io_load(mac_23_26_io_load),
    .io_mulInput(mac_23_26_io_mulInput),
    .io_addInput(mac_23_26_io_addInput),
    .io_output(mac_23_26_io_output),
    .io_passthrough(mac_23_26_io_passthrough)
  );
  MAC mac_23_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_27_clock),
    .reset(mac_23_27_reset),
    .io_load(mac_23_27_io_load),
    .io_mulInput(mac_23_27_io_mulInput),
    .io_addInput(mac_23_27_io_addInput),
    .io_output(mac_23_27_io_output),
    .io_passthrough(mac_23_27_io_passthrough)
  );
  MAC mac_23_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_28_clock),
    .reset(mac_23_28_reset),
    .io_load(mac_23_28_io_load),
    .io_mulInput(mac_23_28_io_mulInput),
    .io_addInput(mac_23_28_io_addInput),
    .io_output(mac_23_28_io_output),
    .io_passthrough(mac_23_28_io_passthrough)
  );
  MAC mac_23_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_29_clock),
    .reset(mac_23_29_reset),
    .io_load(mac_23_29_io_load),
    .io_mulInput(mac_23_29_io_mulInput),
    .io_addInput(mac_23_29_io_addInput),
    .io_output(mac_23_29_io_output),
    .io_passthrough(mac_23_29_io_passthrough)
  );
  MAC mac_23_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_30_clock),
    .reset(mac_23_30_reset),
    .io_load(mac_23_30_io_load),
    .io_mulInput(mac_23_30_io_mulInput),
    .io_addInput(mac_23_30_io_addInput),
    .io_output(mac_23_30_io_output),
    .io_passthrough(mac_23_30_io_passthrough)
  );
  MAC mac_23_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_23_31_clock),
    .reset(mac_23_31_reset),
    .io_load(mac_23_31_io_load),
    .io_mulInput(mac_23_31_io_mulInput),
    .io_addInput(mac_23_31_io_addInput),
    .io_output(mac_23_31_io_output),
    .io_passthrough(mac_23_31_io_passthrough)
  );
  MAC mac_24_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_0_clock),
    .reset(mac_24_0_reset),
    .io_load(mac_24_0_io_load),
    .io_mulInput(mac_24_0_io_mulInput),
    .io_addInput(mac_24_0_io_addInput),
    .io_output(mac_24_0_io_output),
    .io_passthrough(mac_24_0_io_passthrough)
  );
  MAC mac_24_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_1_clock),
    .reset(mac_24_1_reset),
    .io_load(mac_24_1_io_load),
    .io_mulInput(mac_24_1_io_mulInput),
    .io_addInput(mac_24_1_io_addInput),
    .io_output(mac_24_1_io_output),
    .io_passthrough(mac_24_1_io_passthrough)
  );
  MAC mac_24_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_2_clock),
    .reset(mac_24_2_reset),
    .io_load(mac_24_2_io_load),
    .io_mulInput(mac_24_2_io_mulInput),
    .io_addInput(mac_24_2_io_addInput),
    .io_output(mac_24_2_io_output),
    .io_passthrough(mac_24_2_io_passthrough)
  );
  MAC mac_24_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_3_clock),
    .reset(mac_24_3_reset),
    .io_load(mac_24_3_io_load),
    .io_mulInput(mac_24_3_io_mulInput),
    .io_addInput(mac_24_3_io_addInput),
    .io_output(mac_24_3_io_output),
    .io_passthrough(mac_24_3_io_passthrough)
  );
  MAC mac_24_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_4_clock),
    .reset(mac_24_4_reset),
    .io_load(mac_24_4_io_load),
    .io_mulInput(mac_24_4_io_mulInput),
    .io_addInput(mac_24_4_io_addInput),
    .io_output(mac_24_4_io_output),
    .io_passthrough(mac_24_4_io_passthrough)
  );
  MAC mac_24_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_5_clock),
    .reset(mac_24_5_reset),
    .io_load(mac_24_5_io_load),
    .io_mulInput(mac_24_5_io_mulInput),
    .io_addInput(mac_24_5_io_addInput),
    .io_output(mac_24_5_io_output),
    .io_passthrough(mac_24_5_io_passthrough)
  );
  MAC mac_24_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_6_clock),
    .reset(mac_24_6_reset),
    .io_load(mac_24_6_io_load),
    .io_mulInput(mac_24_6_io_mulInput),
    .io_addInput(mac_24_6_io_addInput),
    .io_output(mac_24_6_io_output),
    .io_passthrough(mac_24_6_io_passthrough)
  );
  MAC mac_24_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_7_clock),
    .reset(mac_24_7_reset),
    .io_load(mac_24_7_io_load),
    .io_mulInput(mac_24_7_io_mulInput),
    .io_addInput(mac_24_7_io_addInput),
    .io_output(mac_24_7_io_output),
    .io_passthrough(mac_24_7_io_passthrough)
  );
  MAC mac_24_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_8_clock),
    .reset(mac_24_8_reset),
    .io_load(mac_24_8_io_load),
    .io_mulInput(mac_24_8_io_mulInput),
    .io_addInput(mac_24_8_io_addInput),
    .io_output(mac_24_8_io_output),
    .io_passthrough(mac_24_8_io_passthrough)
  );
  MAC mac_24_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_9_clock),
    .reset(mac_24_9_reset),
    .io_load(mac_24_9_io_load),
    .io_mulInput(mac_24_9_io_mulInput),
    .io_addInput(mac_24_9_io_addInput),
    .io_output(mac_24_9_io_output),
    .io_passthrough(mac_24_9_io_passthrough)
  );
  MAC mac_24_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_10_clock),
    .reset(mac_24_10_reset),
    .io_load(mac_24_10_io_load),
    .io_mulInput(mac_24_10_io_mulInput),
    .io_addInput(mac_24_10_io_addInput),
    .io_output(mac_24_10_io_output),
    .io_passthrough(mac_24_10_io_passthrough)
  );
  MAC mac_24_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_11_clock),
    .reset(mac_24_11_reset),
    .io_load(mac_24_11_io_load),
    .io_mulInput(mac_24_11_io_mulInput),
    .io_addInput(mac_24_11_io_addInput),
    .io_output(mac_24_11_io_output),
    .io_passthrough(mac_24_11_io_passthrough)
  );
  MAC mac_24_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_12_clock),
    .reset(mac_24_12_reset),
    .io_load(mac_24_12_io_load),
    .io_mulInput(mac_24_12_io_mulInput),
    .io_addInput(mac_24_12_io_addInput),
    .io_output(mac_24_12_io_output),
    .io_passthrough(mac_24_12_io_passthrough)
  );
  MAC mac_24_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_13_clock),
    .reset(mac_24_13_reset),
    .io_load(mac_24_13_io_load),
    .io_mulInput(mac_24_13_io_mulInput),
    .io_addInput(mac_24_13_io_addInput),
    .io_output(mac_24_13_io_output),
    .io_passthrough(mac_24_13_io_passthrough)
  );
  MAC mac_24_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_14_clock),
    .reset(mac_24_14_reset),
    .io_load(mac_24_14_io_load),
    .io_mulInput(mac_24_14_io_mulInput),
    .io_addInput(mac_24_14_io_addInput),
    .io_output(mac_24_14_io_output),
    .io_passthrough(mac_24_14_io_passthrough)
  );
  MAC mac_24_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_15_clock),
    .reset(mac_24_15_reset),
    .io_load(mac_24_15_io_load),
    .io_mulInput(mac_24_15_io_mulInput),
    .io_addInput(mac_24_15_io_addInput),
    .io_output(mac_24_15_io_output),
    .io_passthrough(mac_24_15_io_passthrough)
  );
  MAC mac_24_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_16_clock),
    .reset(mac_24_16_reset),
    .io_load(mac_24_16_io_load),
    .io_mulInput(mac_24_16_io_mulInput),
    .io_addInput(mac_24_16_io_addInput),
    .io_output(mac_24_16_io_output),
    .io_passthrough(mac_24_16_io_passthrough)
  );
  MAC mac_24_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_17_clock),
    .reset(mac_24_17_reset),
    .io_load(mac_24_17_io_load),
    .io_mulInput(mac_24_17_io_mulInput),
    .io_addInput(mac_24_17_io_addInput),
    .io_output(mac_24_17_io_output),
    .io_passthrough(mac_24_17_io_passthrough)
  );
  MAC mac_24_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_18_clock),
    .reset(mac_24_18_reset),
    .io_load(mac_24_18_io_load),
    .io_mulInput(mac_24_18_io_mulInput),
    .io_addInput(mac_24_18_io_addInput),
    .io_output(mac_24_18_io_output),
    .io_passthrough(mac_24_18_io_passthrough)
  );
  MAC mac_24_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_19_clock),
    .reset(mac_24_19_reset),
    .io_load(mac_24_19_io_load),
    .io_mulInput(mac_24_19_io_mulInput),
    .io_addInput(mac_24_19_io_addInput),
    .io_output(mac_24_19_io_output),
    .io_passthrough(mac_24_19_io_passthrough)
  );
  MAC mac_24_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_20_clock),
    .reset(mac_24_20_reset),
    .io_load(mac_24_20_io_load),
    .io_mulInput(mac_24_20_io_mulInput),
    .io_addInput(mac_24_20_io_addInput),
    .io_output(mac_24_20_io_output),
    .io_passthrough(mac_24_20_io_passthrough)
  );
  MAC mac_24_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_21_clock),
    .reset(mac_24_21_reset),
    .io_load(mac_24_21_io_load),
    .io_mulInput(mac_24_21_io_mulInput),
    .io_addInput(mac_24_21_io_addInput),
    .io_output(mac_24_21_io_output),
    .io_passthrough(mac_24_21_io_passthrough)
  );
  MAC mac_24_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_22_clock),
    .reset(mac_24_22_reset),
    .io_load(mac_24_22_io_load),
    .io_mulInput(mac_24_22_io_mulInput),
    .io_addInput(mac_24_22_io_addInput),
    .io_output(mac_24_22_io_output),
    .io_passthrough(mac_24_22_io_passthrough)
  );
  MAC mac_24_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_23_clock),
    .reset(mac_24_23_reset),
    .io_load(mac_24_23_io_load),
    .io_mulInput(mac_24_23_io_mulInput),
    .io_addInput(mac_24_23_io_addInput),
    .io_output(mac_24_23_io_output),
    .io_passthrough(mac_24_23_io_passthrough)
  );
  MAC mac_24_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_24_clock),
    .reset(mac_24_24_reset),
    .io_load(mac_24_24_io_load),
    .io_mulInput(mac_24_24_io_mulInput),
    .io_addInput(mac_24_24_io_addInput),
    .io_output(mac_24_24_io_output),
    .io_passthrough(mac_24_24_io_passthrough)
  );
  MAC mac_24_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_25_clock),
    .reset(mac_24_25_reset),
    .io_load(mac_24_25_io_load),
    .io_mulInput(mac_24_25_io_mulInput),
    .io_addInput(mac_24_25_io_addInput),
    .io_output(mac_24_25_io_output),
    .io_passthrough(mac_24_25_io_passthrough)
  );
  MAC mac_24_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_26_clock),
    .reset(mac_24_26_reset),
    .io_load(mac_24_26_io_load),
    .io_mulInput(mac_24_26_io_mulInput),
    .io_addInput(mac_24_26_io_addInput),
    .io_output(mac_24_26_io_output),
    .io_passthrough(mac_24_26_io_passthrough)
  );
  MAC mac_24_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_27_clock),
    .reset(mac_24_27_reset),
    .io_load(mac_24_27_io_load),
    .io_mulInput(mac_24_27_io_mulInput),
    .io_addInput(mac_24_27_io_addInput),
    .io_output(mac_24_27_io_output),
    .io_passthrough(mac_24_27_io_passthrough)
  );
  MAC mac_24_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_28_clock),
    .reset(mac_24_28_reset),
    .io_load(mac_24_28_io_load),
    .io_mulInput(mac_24_28_io_mulInput),
    .io_addInput(mac_24_28_io_addInput),
    .io_output(mac_24_28_io_output),
    .io_passthrough(mac_24_28_io_passthrough)
  );
  MAC mac_24_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_29_clock),
    .reset(mac_24_29_reset),
    .io_load(mac_24_29_io_load),
    .io_mulInput(mac_24_29_io_mulInput),
    .io_addInput(mac_24_29_io_addInput),
    .io_output(mac_24_29_io_output),
    .io_passthrough(mac_24_29_io_passthrough)
  );
  MAC mac_24_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_30_clock),
    .reset(mac_24_30_reset),
    .io_load(mac_24_30_io_load),
    .io_mulInput(mac_24_30_io_mulInput),
    .io_addInput(mac_24_30_io_addInput),
    .io_output(mac_24_30_io_output),
    .io_passthrough(mac_24_30_io_passthrough)
  );
  MAC mac_24_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_24_31_clock),
    .reset(mac_24_31_reset),
    .io_load(mac_24_31_io_load),
    .io_mulInput(mac_24_31_io_mulInput),
    .io_addInput(mac_24_31_io_addInput),
    .io_output(mac_24_31_io_output),
    .io_passthrough(mac_24_31_io_passthrough)
  );
  MAC mac_25_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_0_clock),
    .reset(mac_25_0_reset),
    .io_load(mac_25_0_io_load),
    .io_mulInput(mac_25_0_io_mulInput),
    .io_addInput(mac_25_0_io_addInput),
    .io_output(mac_25_0_io_output),
    .io_passthrough(mac_25_0_io_passthrough)
  );
  MAC mac_25_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_1_clock),
    .reset(mac_25_1_reset),
    .io_load(mac_25_1_io_load),
    .io_mulInput(mac_25_1_io_mulInput),
    .io_addInput(mac_25_1_io_addInput),
    .io_output(mac_25_1_io_output),
    .io_passthrough(mac_25_1_io_passthrough)
  );
  MAC mac_25_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_2_clock),
    .reset(mac_25_2_reset),
    .io_load(mac_25_2_io_load),
    .io_mulInput(mac_25_2_io_mulInput),
    .io_addInput(mac_25_2_io_addInput),
    .io_output(mac_25_2_io_output),
    .io_passthrough(mac_25_2_io_passthrough)
  );
  MAC mac_25_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_3_clock),
    .reset(mac_25_3_reset),
    .io_load(mac_25_3_io_load),
    .io_mulInput(mac_25_3_io_mulInput),
    .io_addInput(mac_25_3_io_addInput),
    .io_output(mac_25_3_io_output),
    .io_passthrough(mac_25_3_io_passthrough)
  );
  MAC mac_25_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_4_clock),
    .reset(mac_25_4_reset),
    .io_load(mac_25_4_io_load),
    .io_mulInput(mac_25_4_io_mulInput),
    .io_addInput(mac_25_4_io_addInput),
    .io_output(mac_25_4_io_output),
    .io_passthrough(mac_25_4_io_passthrough)
  );
  MAC mac_25_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_5_clock),
    .reset(mac_25_5_reset),
    .io_load(mac_25_5_io_load),
    .io_mulInput(mac_25_5_io_mulInput),
    .io_addInput(mac_25_5_io_addInput),
    .io_output(mac_25_5_io_output),
    .io_passthrough(mac_25_5_io_passthrough)
  );
  MAC mac_25_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_6_clock),
    .reset(mac_25_6_reset),
    .io_load(mac_25_6_io_load),
    .io_mulInput(mac_25_6_io_mulInput),
    .io_addInput(mac_25_6_io_addInput),
    .io_output(mac_25_6_io_output),
    .io_passthrough(mac_25_6_io_passthrough)
  );
  MAC mac_25_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_7_clock),
    .reset(mac_25_7_reset),
    .io_load(mac_25_7_io_load),
    .io_mulInput(mac_25_7_io_mulInput),
    .io_addInput(mac_25_7_io_addInput),
    .io_output(mac_25_7_io_output),
    .io_passthrough(mac_25_7_io_passthrough)
  );
  MAC mac_25_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_8_clock),
    .reset(mac_25_8_reset),
    .io_load(mac_25_8_io_load),
    .io_mulInput(mac_25_8_io_mulInput),
    .io_addInput(mac_25_8_io_addInput),
    .io_output(mac_25_8_io_output),
    .io_passthrough(mac_25_8_io_passthrough)
  );
  MAC mac_25_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_9_clock),
    .reset(mac_25_9_reset),
    .io_load(mac_25_9_io_load),
    .io_mulInput(mac_25_9_io_mulInput),
    .io_addInput(mac_25_9_io_addInput),
    .io_output(mac_25_9_io_output),
    .io_passthrough(mac_25_9_io_passthrough)
  );
  MAC mac_25_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_10_clock),
    .reset(mac_25_10_reset),
    .io_load(mac_25_10_io_load),
    .io_mulInput(mac_25_10_io_mulInput),
    .io_addInput(mac_25_10_io_addInput),
    .io_output(mac_25_10_io_output),
    .io_passthrough(mac_25_10_io_passthrough)
  );
  MAC mac_25_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_11_clock),
    .reset(mac_25_11_reset),
    .io_load(mac_25_11_io_load),
    .io_mulInput(mac_25_11_io_mulInput),
    .io_addInput(mac_25_11_io_addInput),
    .io_output(mac_25_11_io_output),
    .io_passthrough(mac_25_11_io_passthrough)
  );
  MAC mac_25_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_12_clock),
    .reset(mac_25_12_reset),
    .io_load(mac_25_12_io_load),
    .io_mulInput(mac_25_12_io_mulInput),
    .io_addInput(mac_25_12_io_addInput),
    .io_output(mac_25_12_io_output),
    .io_passthrough(mac_25_12_io_passthrough)
  );
  MAC mac_25_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_13_clock),
    .reset(mac_25_13_reset),
    .io_load(mac_25_13_io_load),
    .io_mulInput(mac_25_13_io_mulInput),
    .io_addInput(mac_25_13_io_addInput),
    .io_output(mac_25_13_io_output),
    .io_passthrough(mac_25_13_io_passthrough)
  );
  MAC mac_25_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_14_clock),
    .reset(mac_25_14_reset),
    .io_load(mac_25_14_io_load),
    .io_mulInput(mac_25_14_io_mulInput),
    .io_addInput(mac_25_14_io_addInput),
    .io_output(mac_25_14_io_output),
    .io_passthrough(mac_25_14_io_passthrough)
  );
  MAC mac_25_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_15_clock),
    .reset(mac_25_15_reset),
    .io_load(mac_25_15_io_load),
    .io_mulInput(mac_25_15_io_mulInput),
    .io_addInput(mac_25_15_io_addInput),
    .io_output(mac_25_15_io_output),
    .io_passthrough(mac_25_15_io_passthrough)
  );
  MAC mac_25_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_16_clock),
    .reset(mac_25_16_reset),
    .io_load(mac_25_16_io_load),
    .io_mulInput(mac_25_16_io_mulInput),
    .io_addInput(mac_25_16_io_addInput),
    .io_output(mac_25_16_io_output),
    .io_passthrough(mac_25_16_io_passthrough)
  );
  MAC mac_25_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_17_clock),
    .reset(mac_25_17_reset),
    .io_load(mac_25_17_io_load),
    .io_mulInput(mac_25_17_io_mulInput),
    .io_addInput(mac_25_17_io_addInput),
    .io_output(mac_25_17_io_output),
    .io_passthrough(mac_25_17_io_passthrough)
  );
  MAC mac_25_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_18_clock),
    .reset(mac_25_18_reset),
    .io_load(mac_25_18_io_load),
    .io_mulInput(mac_25_18_io_mulInput),
    .io_addInput(mac_25_18_io_addInput),
    .io_output(mac_25_18_io_output),
    .io_passthrough(mac_25_18_io_passthrough)
  );
  MAC mac_25_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_19_clock),
    .reset(mac_25_19_reset),
    .io_load(mac_25_19_io_load),
    .io_mulInput(mac_25_19_io_mulInput),
    .io_addInput(mac_25_19_io_addInput),
    .io_output(mac_25_19_io_output),
    .io_passthrough(mac_25_19_io_passthrough)
  );
  MAC mac_25_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_20_clock),
    .reset(mac_25_20_reset),
    .io_load(mac_25_20_io_load),
    .io_mulInput(mac_25_20_io_mulInput),
    .io_addInput(mac_25_20_io_addInput),
    .io_output(mac_25_20_io_output),
    .io_passthrough(mac_25_20_io_passthrough)
  );
  MAC mac_25_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_21_clock),
    .reset(mac_25_21_reset),
    .io_load(mac_25_21_io_load),
    .io_mulInput(mac_25_21_io_mulInput),
    .io_addInput(mac_25_21_io_addInput),
    .io_output(mac_25_21_io_output),
    .io_passthrough(mac_25_21_io_passthrough)
  );
  MAC mac_25_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_22_clock),
    .reset(mac_25_22_reset),
    .io_load(mac_25_22_io_load),
    .io_mulInput(mac_25_22_io_mulInput),
    .io_addInput(mac_25_22_io_addInput),
    .io_output(mac_25_22_io_output),
    .io_passthrough(mac_25_22_io_passthrough)
  );
  MAC mac_25_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_23_clock),
    .reset(mac_25_23_reset),
    .io_load(mac_25_23_io_load),
    .io_mulInput(mac_25_23_io_mulInput),
    .io_addInput(mac_25_23_io_addInput),
    .io_output(mac_25_23_io_output),
    .io_passthrough(mac_25_23_io_passthrough)
  );
  MAC mac_25_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_24_clock),
    .reset(mac_25_24_reset),
    .io_load(mac_25_24_io_load),
    .io_mulInput(mac_25_24_io_mulInput),
    .io_addInput(mac_25_24_io_addInput),
    .io_output(mac_25_24_io_output),
    .io_passthrough(mac_25_24_io_passthrough)
  );
  MAC mac_25_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_25_clock),
    .reset(mac_25_25_reset),
    .io_load(mac_25_25_io_load),
    .io_mulInput(mac_25_25_io_mulInput),
    .io_addInput(mac_25_25_io_addInput),
    .io_output(mac_25_25_io_output),
    .io_passthrough(mac_25_25_io_passthrough)
  );
  MAC mac_25_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_26_clock),
    .reset(mac_25_26_reset),
    .io_load(mac_25_26_io_load),
    .io_mulInput(mac_25_26_io_mulInput),
    .io_addInput(mac_25_26_io_addInput),
    .io_output(mac_25_26_io_output),
    .io_passthrough(mac_25_26_io_passthrough)
  );
  MAC mac_25_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_27_clock),
    .reset(mac_25_27_reset),
    .io_load(mac_25_27_io_load),
    .io_mulInput(mac_25_27_io_mulInput),
    .io_addInput(mac_25_27_io_addInput),
    .io_output(mac_25_27_io_output),
    .io_passthrough(mac_25_27_io_passthrough)
  );
  MAC mac_25_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_28_clock),
    .reset(mac_25_28_reset),
    .io_load(mac_25_28_io_load),
    .io_mulInput(mac_25_28_io_mulInput),
    .io_addInput(mac_25_28_io_addInput),
    .io_output(mac_25_28_io_output),
    .io_passthrough(mac_25_28_io_passthrough)
  );
  MAC mac_25_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_29_clock),
    .reset(mac_25_29_reset),
    .io_load(mac_25_29_io_load),
    .io_mulInput(mac_25_29_io_mulInput),
    .io_addInput(mac_25_29_io_addInput),
    .io_output(mac_25_29_io_output),
    .io_passthrough(mac_25_29_io_passthrough)
  );
  MAC mac_25_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_30_clock),
    .reset(mac_25_30_reset),
    .io_load(mac_25_30_io_load),
    .io_mulInput(mac_25_30_io_mulInput),
    .io_addInput(mac_25_30_io_addInput),
    .io_output(mac_25_30_io_output),
    .io_passthrough(mac_25_30_io_passthrough)
  );
  MAC mac_25_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_25_31_clock),
    .reset(mac_25_31_reset),
    .io_load(mac_25_31_io_load),
    .io_mulInput(mac_25_31_io_mulInput),
    .io_addInput(mac_25_31_io_addInput),
    .io_output(mac_25_31_io_output),
    .io_passthrough(mac_25_31_io_passthrough)
  );
  MAC mac_26_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_0_clock),
    .reset(mac_26_0_reset),
    .io_load(mac_26_0_io_load),
    .io_mulInput(mac_26_0_io_mulInput),
    .io_addInput(mac_26_0_io_addInput),
    .io_output(mac_26_0_io_output),
    .io_passthrough(mac_26_0_io_passthrough)
  );
  MAC mac_26_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_1_clock),
    .reset(mac_26_1_reset),
    .io_load(mac_26_1_io_load),
    .io_mulInput(mac_26_1_io_mulInput),
    .io_addInput(mac_26_1_io_addInput),
    .io_output(mac_26_1_io_output),
    .io_passthrough(mac_26_1_io_passthrough)
  );
  MAC mac_26_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_2_clock),
    .reset(mac_26_2_reset),
    .io_load(mac_26_2_io_load),
    .io_mulInput(mac_26_2_io_mulInput),
    .io_addInput(mac_26_2_io_addInput),
    .io_output(mac_26_2_io_output),
    .io_passthrough(mac_26_2_io_passthrough)
  );
  MAC mac_26_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_3_clock),
    .reset(mac_26_3_reset),
    .io_load(mac_26_3_io_load),
    .io_mulInput(mac_26_3_io_mulInput),
    .io_addInput(mac_26_3_io_addInput),
    .io_output(mac_26_3_io_output),
    .io_passthrough(mac_26_3_io_passthrough)
  );
  MAC mac_26_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_4_clock),
    .reset(mac_26_4_reset),
    .io_load(mac_26_4_io_load),
    .io_mulInput(mac_26_4_io_mulInput),
    .io_addInput(mac_26_4_io_addInput),
    .io_output(mac_26_4_io_output),
    .io_passthrough(mac_26_4_io_passthrough)
  );
  MAC mac_26_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_5_clock),
    .reset(mac_26_5_reset),
    .io_load(mac_26_5_io_load),
    .io_mulInput(mac_26_5_io_mulInput),
    .io_addInput(mac_26_5_io_addInput),
    .io_output(mac_26_5_io_output),
    .io_passthrough(mac_26_5_io_passthrough)
  );
  MAC mac_26_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_6_clock),
    .reset(mac_26_6_reset),
    .io_load(mac_26_6_io_load),
    .io_mulInput(mac_26_6_io_mulInput),
    .io_addInput(mac_26_6_io_addInput),
    .io_output(mac_26_6_io_output),
    .io_passthrough(mac_26_6_io_passthrough)
  );
  MAC mac_26_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_7_clock),
    .reset(mac_26_7_reset),
    .io_load(mac_26_7_io_load),
    .io_mulInput(mac_26_7_io_mulInput),
    .io_addInput(mac_26_7_io_addInput),
    .io_output(mac_26_7_io_output),
    .io_passthrough(mac_26_7_io_passthrough)
  );
  MAC mac_26_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_8_clock),
    .reset(mac_26_8_reset),
    .io_load(mac_26_8_io_load),
    .io_mulInput(mac_26_8_io_mulInput),
    .io_addInput(mac_26_8_io_addInput),
    .io_output(mac_26_8_io_output),
    .io_passthrough(mac_26_8_io_passthrough)
  );
  MAC mac_26_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_9_clock),
    .reset(mac_26_9_reset),
    .io_load(mac_26_9_io_load),
    .io_mulInput(mac_26_9_io_mulInput),
    .io_addInput(mac_26_9_io_addInput),
    .io_output(mac_26_9_io_output),
    .io_passthrough(mac_26_9_io_passthrough)
  );
  MAC mac_26_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_10_clock),
    .reset(mac_26_10_reset),
    .io_load(mac_26_10_io_load),
    .io_mulInput(mac_26_10_io_mulInput),
    .io_addInput(mac_26_10_io_addInput),
    .io_output(mac_26_10_io_output),
    .io_passthrough(mac_26_10_io_passthrough)
  );
  MAC mac_26_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_11_clock),
    .reset(mac_26_11_reset),
    .io_load(mac_26_11_io_load),
    .io_mulInput(mac_26_11_io_mulInput),
    .io_addInput(mac_26_11_io_addInput),
    .io_output(mac_26_11_io_output),
    .io_passthrough(mac_26_11_io_passthrough)
  );
  MAC mac_26_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_12_clock),
    .reset(mac_26_12_reset),
    .io_load(mac_26_12_io_load),
    .io_mulInput(mac_26_12_io_mulInput),
    .io_addInput(mac_26_12_io_addInput),
    .io_output(mac_26_12_io_output),
    .io_passthrough(mac_26_12_io_passthrough)
  );
  MAC mac_26_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_13_clock),
    .reset(mac_26_13_reset),
    .io_load(mac_26_13_io_load),
    .io_mulInput(mac_26_13_io_mulInput),
    .io_addInput(mac_26_13_io_addInput),
    .io_output(mac_26_13_io_output),
    .io_passthrough(mac_26_13_io_passthrough)
  );
  MAC mac_26_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_14_clock),
    .reset(mac_26_14_reset),
    .io_load(mac_26_14_io_load),
    .io_mulInput(mac_26_14_io_mulInput),
    .io_addInput(mac_26_14_io_addInput),
    .io_output(mac_26_14_io_output),
    .io_passthrough(mac_26_14_io_passthrough)
  );
  MAC mac_26_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_15_clock),
    .reset(mac_26_15_reset),
    .io_load(mac_26_15_io_load),
    .io_mulInput(mac_26_15_io_mulInput),
    .io_addInput(mac_26_15_io_addInput),
    .io_output(mac_26_15_io_output),
    .io_passthrough(mac_26_15_io_passthrough)
  );
  MAC mac_26_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_16_clock),
    .reset(mac_26_16_reset),
    .io_load(mac_26_16_io_load),
    .io_mulInput(mac_26_16_io_mulInput),
    .io_addInput(mac_26_16_io_addInput),
    .io_output(mac_26_16_io_output),
    .io_passthrough(mac_26_16_io_passthrough)
  );
  MAC mac_26_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_17_clock),
    .reset(mac_26_17_reset),
    .io_load(mac_26_17_io_load),
    .io_mulInput(mac_26_17_io_mulInput),
    .io_addInput(mac_26_17_io_addInput),
    .io_output(mac_26_17_io_output),
    .io_passthrough(mac_26_17_io_passthrough)
  );
  MAC mac_26_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_18_clock),
    .reset(mac_26_18_reset),
    .io_load(mac_26_18_io_load),
    .io_mulInput(mac_26_18_io_mulInput),
    .io_addInput(mac_26_18_io_addInput),
    .io_output(mac_26_18_io_output),
    .io_passthrough(mac_26_18_io_passthrough)
  );
  MAC mac_26_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_19_clock),
    .reset(mac_26_19_reset),
    .io_load(mac_26_19_io_load),
    .io_mulInput(mac_26_19_io_mulInput),
    .io_addInput(mac_26_19_io_addInput),
    .io_output(mac_26_19_io_output),
    .io_passthrough(mac_26_19_io_passthrough)
  );
  MAC mac_26_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_20_clock),
    .reset(mac_26_20_reset),
    .io_load(mac_26_20_io_load),
    .io_mulInput(mac_26_20_io_mulInput),
    .io_addInput(mac_26_20_io_addInput),
    .io_output(mac_26_20_io_output),
    .io_passthrough(mac_26_20_io_passthrough)
  );
  MAC mac_26_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_21_clock),
    .reset(mac_26_21_reset),
    .io_load(mac_26_21_io_load),
    .io_mulInput(mac_26_21_io_mulInput),
    .io_addInput(mac_26_21_io_addInput),
    .io_output(mac_26_21_io_output),
    .io_passthrough(mac_26_21_io_passthrough)
  );
  MAC mac_26_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_22_clock),
    .reset(mac_26_22_reset),
    .io_load(mac_26_22_io_load),
    .io_mulInput(mac_26_22_io_mulInput),
    .io_addInput(mac_26_22_io_addInput),
    .io_output(mac_26_22_io_output),
    .io_passthrough(mac_26_22_io_passthrough)
  );
  MAC mac_26_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_23_clock),
    .reset(mac_26_23_reset),
    .io_load(mac_26_23_io_load),
    .io_mulInput(mac_26_23_io_mulInput),
    .io_addInput(mac_26_23_io_addInput),
    .io_output(mac_26_23_io_output),
    .io_passthrough(mac_26_23_io_passthrough)
  );
  MAC mac_26_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_24_clock),
    .reset(mac_26_24_reset),
    .io_load(mac_26_24_io_load),
    .io_mulInput(mac_26_24_io_mulInput),
    .io_addInput(mac_26_24_io_addInput),
    .io_output(mac_26_24_io_output),
    .io_passthrough(mac_26_24_io_passthrough)
  );
  MAC mac_26_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_25_clock),
    .reset(mac_26_25_reset),
    .io_load(mac_26_25_io_load),
    .io_mulInput(mac_26_25_io_mulInput),
    .io_addInput(mac_26_25_io_addInput),
    .io_output(mac_26_25_io_output),
    .io_passthrough(mac_26_25_io_passthrough)
  );
  MAC mac_26_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_26_clock),
    .reset(mac_26_26_reset),
    .io_load(mac_26_26_io_load),
    .io_mulInput(mac_26_26_io_mulInput),
    .io_addInput(mac_26_26_io_addInput),
    .io_output(mac_26_26_io_output),
    .io_passthrough(mac_26_26_io_passthrough)
  );
  MAC mac_26_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_27_clock),
    .reset(mac_26_27_reset),
    .io_load(mac_26_27_io_load),
    .io_mulInput(mac_26_27_io_mulInput),
    .io_addInput(mac_26_27_io_addInput),
    .io_output(mac_26_27_io_output),
    .io_passthrough(mac_26_27_io_passthrough)
  );
  MAC mac_26_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_28_clock),
    .reset(mac_26_28_reset),
    .io_load(mac_26_28_io_load),
    .io_mulInput(mac_26_28_io_mulInput),
    .io_addInput(mac_26_28_io_addInput),
    .io_output(mac_26_28_io_output),
    .io_passthrough(mac_26_28_io_passthrough)
  );
  MAC mac_26_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_29_clock),
    .reset(mac_26_29_reset),
    .io_load(mac_26_29_io_load),
    .io_mulInput(mac_26_29_io_mulInput),
    .io_addInput(mac_26_29_io_addInput),
    .io_output(mac_26_29_io_output),
    .io_passthrough(mac_26_29_io_passthrough)
  );
  MAC mac_26_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_30_clock),
    .reset(mac_26_30_reset),
    .io_load(mac_26_30_io_load),
    .io_mulInput(mac_26_30_io_mulInput),
    .io_addInput(mac_26_30_io_addInput),
    .io_output(mac_26_30_io_output),
    .io_passthrough(mac_26_30_io_passthrough)
  );
  MAC mac_26_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_26_31_clock),
    .reset(mac_26_31_reset),
    .io_load(mac_26_31_io_load),
    .io_mulInput(mac_26_31_io_mulInput),
    .io_addInput(mac_26_31_io_addInput),
    .io_output(mac_26_31_io_output),
    .io_passthrough(mac_26_31_io_passthrough)
  );
  MAC mac_27_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_0_clock),
    .reset(mac_27_0_reset),
    .io_load(mac_27_0_io_load),
    .io_mulInput(mac_27_0_io_mulInput),
    .io_addInput(mac_27_0_io_addInput),
    .io_output(mac_27_0_io_output),
    .io_passthrough(mac_27_0_io_passthrough)
  );
  MAC mac_27_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_1_clock),
    .reset(mac_27_1_reset),
    .io_load(mac_27_1_io_load),
    .io_mulInput(mac_27_1_io_mulInput),
    .io_addInput(mac_27_1_io_addInput),
    .io_output(mac_27_1_io_output),
    .io_passthrough(mac_27_1_io_passthrough)
  );
  MAC mac_27_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_2_clock),
    .reset(mac_27_2_reset),
    .io_load(mac_27_2_io_load),
    .io_mulInput(mac_27_2_io_mulInput),
    .io_addInput(mac_27_2_io_addInput),
    .io_output(mac_27_2_io_output),
    .io_passthrough(mac_27_2_io_passthrough)
  );
  MAC mac_27_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_3_clock),
    .reset(mac_27_3_reset),
    .io_load(mac_27_3_io_load),
    .io_mulInput(mac_27_3_io_mulInput),
    .io_addInput(mac_27_3_io_addInput),
    .io_output(mac_27_3_io_output),
    .io_passthrough(mac_27_3_io_passthrough)
  );
  MAC mac_27_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_4_clock),
    .reset(mac_27_4_reset),
    .io_load(mac_27_4_io_load),
    .io_mulInput(mac_27_4_io_mulInput),
    .io_addInput(mac_27_4_io_addInput),
    .io_output(mac_27_4_io_output),
    .io_passthrough(mac_27_4_io_passthrough)
  );
  MAC mac_27_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_5_clock),
    .reset(mac_27_5_reset),
    .io_load(mac_27_5_io_load),
    .io_mulInput(mac_27_5_io_mulInput),
    .io_addInput(mac_27_5_io_addInput),
    .io_output(mac_27_5_io_output),
    .io_passthrough(mac_27_5_io_passthrough)
  );
  MAC mac_27_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_6_clock),
    .reset(mac_27_6_reset),
    .io_load(mac_27_6_io_load),
    .io_mulInput(mac_27_6_io_mulInput),
    .io_addInput(mac_27_6_io_addInput),
    .io_output(mac_27_6_io_output),
    .io_passthrough(mac_27_6_io_passthrough)
  );
  MAC mac_27_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_7_clock),
    .reset(mac_27_7_reset),
    .io_load(mac_27_7_io_load),
    .io_mulInput(mac_27_7_io_mulInput),
    .io_addInput(mac_27_7_io_addInput),
    .io_output(mac_27_7_io_output),
    .io_passthrough(mac_27_7_io_passthrough)
  );
  MAC mac_27_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_8_clock),
    .reset(mac_27_8_reset),
    .io_load(mac_27_8_io_load),
    .io_mulInput(mac_27_8_io_mulInput),
    .io_addInput(mac_27_8_io_addInput),
    .io_output(mac_27_8_io_output),
    .io_passthrough(mac_27_8_io_passthrough)
  );
  MAC mac_27_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_9_clock),
    .reset(mac_27_9_reset),
    .io_load(mac_27_9_io_load),
    .io_mulInput(mac_27_9_io_mulInput),
    .io_addInput(mac_27_9_io_addInput),
    .io_output(mac_27_9_io_output),
    .io_passthrough(mac_27_9_io_passthrough)
  );
  MAC mac_27_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_10_clock),
    .reset(mac_27_10_reset),
    .io_load(mac_27_10_io_load),
    .io_mulInput(mac_27_10_io_mulInput),
    .io_addInput(mac_27_10_io_addInput),
    .io_output(mac_27_10_io_output),
    .io_passthrough(mac_27_10_io_passthrough)
  );
  MAC mac_27_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_11_clock),
    .reset(mac_27_11_reset),
    .io_load(mac_27_11_io_load),
    .io_mulInput(mac_27_11_io_mulInput),
    .io_addInput(mac_27_11_io_addInput),
    .io_output(mac_27_11_io_output),
    .io_passthrough(mac_27_11_io_passthrough)
  );
  MAC mac_27_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_12_clock),
    .reset(mac_27_12_reset),
    .io_load(mac_27_12_io_load),
    .io_mulInput(mac_27_12_io_mulInput),
    .io_addInput(mac_27_12_io_addInput),
    .io_output(mac_27_12_io_output),
    .io_passthrough(mac_27_12_io_passthrough)
  );
  MAC mac_27_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_13_clock),
    .reset(mac_27_13_reset),
    .io_load(mac_27_13_io_load),
    .io_mulInput(mac_27_13_io_mulInput),
    .io_addInput(mac_27_13_io_addInput),
    .io_output(mac_27_13_io_output),
    .io_passthrough(mac_27_13_io_passthrough)
  );
  MAC mac_27_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_14_clock),
    .reset(mac_27_14_reset),
    .io_load(mac_27_14_io_load),
    .io_mulInput(mac_27_14_io_mulInput),
    .io_addInput(mac_27_14_io_addInput),
    .io_output(mac_27_14_io_output),
    .io_passthrough(mac_27_14_io_passthrough)
  );
  MAC mac_27_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_15_clock),
    .reset(mac_27_15_reset),
    .io_load(mac_27_15_io_load),
    .io_mulInput(mac_27_15_io_mulInput),
    .io_addInput(mac_27_15_io_addInput),
    .io_output(mac_27_15_io_output),
    .io_passthrough(mac_27_15_io_passthrough)
  );
  MAC mac_27_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_16_clock),
    .reset(mac_27_16_reset),
    .io_load(mac_27_16_io_load),
    .io_mulInput(mac_27_16_io_mulInput),
    .io_addInput(mac_27_16_io_addInput),
    .io_output(mac_27_16_io_output),
    .io_passthrough(mac_27_16_io_passthrough)
  );
  MAC mac_27_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_17_clock),
    .reset(mac_27_17_reset),
    .io_load(mac_27_17_io_load),
    .io_mulInput(mac_27_17_io_mulInput),
    .io_addInput(mac_27_17_io_addInput),
    .io_output(mac_27_17_io_output),
    .io_passthrough(mac_27_17_io_passthrough)
  );
  MAC mac_27_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_18_clock),
    .reset(mac_27_18_reset),
    .io_load(mac_27_18_io_load),
    .io_mulInput(mac_27_18_io_mulInput),
    .io_addInput(mac_27_18_io_addInput),
    .io_output(mac_27_18_io_output),
    .io_passthrough(mac_27_18_io_passthrough)
  );
  MAC mac_27_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_19_clock),
    .reset(mac_27_19_reset),
    .io_load(mac_27_19_io_load),
    .io_mulInput(mac_27_19_io_mulInput),
    .io_addInput(mac_27_19_io_addInput),
    .io_output(mac_27_19_io_output),
    .io_passthrough(mac_27_19_io_passthrough)
  );
  MAC mac_27_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_20_clock),
    .reset(mac_27_20_reset),
    .io_load(mac_27_20_io_load),
    .io_mulInput(mac_27_20_io_mulInput),
    .io_addInput(mac_27_20_io_addInput),
    .io_output(mac_27_20_io_output),
    .io_passthrough(mac_27_20_io_passthrough)
  );
  MAC mac_27_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_21_clock),
    .reset(mac_27_21_reset),
    .io_load(mac_27_21_io_load),
    .io_mulInput(mac_27_21_io_mulInput),
    .io_addInput(mac_27_21_io_addInput),
    .io_output(mac_27_21_io_output),
    .io_passthrough(mac_27_21_io_passthrough)
  );
  MAC mac_27_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_22_clock),
    .reset(mac_27_22_reset),
    .io_load(mac_27_22_io_load),
    .io_mulInput(mac_27_22_io_mulInput),
    .io_addInput(mac_27_22_io_addInput),
    .io_output(mac_27_22_io_output),
    .io_passthrough(mac_27_22_io_passthrough)
  );
  MAC mac_27_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_23_clock),
    .reset(mac_27_23_reset),
    .io_load(mac_27_23_io_load),
    .io_mulInput(mac_27_23_io_mulInput),
    .io_addInput(mac_27_23_io_addInput),
    .io_output(mac_27_23_io_output),
    .io_passthrough(mac_27_23_io_passthrough)
  );
  MAC mac_27_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_24_clock),
    .reset(mac_27_24_reset),
    .io_load(mac_27_24_io_load),
    .io_mulInput(mac_27_24_io_mulInput),
    .io_addInput(mac_27_24_io_addInput),
    .io_output(mac_27_24_io_output),
    .io_passthrough(mac_27_24_io_passthrough)
  );
  MAC mac_27_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_25_clock),
    .reset(mac_27_25_reset),
    .io_load(mac_27_25_io_load),
    .io_mulInput(mac_27_25_io_mulInput),
    .io_addInput(mac_27_25_io_addInput),
    .io_output(mac_27_25_io_output),
    .io_passthrough(mac_27_25_io_passthrough)
  );
  MAC mac_27_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_26_clock),
    .reset(mac_27_26_reset),
    .io_load(mac_27_26_io_load),
    .io_mulInput(mac_27_26_io_mulInput),
    .io_addInput(mac_27_26_io_addInput),
    .io_output(mac_27_26_io_output),
    .io_passthrough(mac_27_26_io_passthrough)
  );
  MAC mac_27_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_27_clock),
    .reset(mac_27_27_reset),
    .io_load(mac_27_27_io_load),
    .io_mulInput(mac_27_27_io_mulInput),
    .io_addInput(mac_27_27_io_addInput),
    .io_output(mac_27_27_io_output),
    .io_passthrough(mac_27_27_io_passthrough)
  );
  MAC mac_27_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_28_clock),
    .reset(mac_27_28_reset),
    .io_load(mac_27_28_io_load),
    .io_mulInput(mac_27_28_io_mulInput),
    .io_addInput(mac_27_28_io_addInput),
    .io_output(mac_27_28_io_output),
    .io_passthrough(mac_27_28_io_passthrough)
  );
  MAC mac_27_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_29_clock),
    .reset(mac_27_29_reset),
    .io_load(mac_27_29_io_load),
    .io_mulInput(mac_27_29_io_mulInput),
    .io_addInput(mac_27_29_io_addInput),
    .io_output(mac_27_29_io_output),
    .io_passthrough(mac_27_29_io_passthrough)
  );
  MAC mac_27_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_30_clock),
    .reset(mac_27_30_reset),
    .io_load(mac_27_30_io_load),
    .io_mulInput(mac_27_30_io_mulInput),
    .io_addInput(mac_27_30_io_addInput),
    .io_output(mac_27_30_io_output),
    .io_passthrough(mac_27_30_io_passthrough)
  );
  MAC mac_27_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_27_31_clock),
    .reset(mac_27_31_reset),
    .io_load(mac_27_31_io_load),
    .io_mulInput(mac_27_31_io_mulInput),
    .io_addInput(mac_27_31_io_addInput),
    .io_output(mac_27_31_io_output),
    .io_passthrough(mac_27_31_io_passthrough)
  );
  MAC mac_28_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_0_clock),
    .reset(mac_28_0_reset),
    .io_load(mac_28_0_io_load),
    .io_mulInput(mac_28_0_io_mulInput),
    .io_addInput(mac_28_0_io_addInput),
    .io_output(mac_28_0_io_output),
    .io_passthrough(mac_28_0_io_passthrough)
  );
  MAC mac_28_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_1_clock),
    .reset(mac_28_1_reset),
    .io_load(mac_28_1_io_load),
    .io_mulInput(mac_28_1_io_mulInput),
    .io_addInput(mac_28_1_io_addInput),
    .io_output(mac_28_1_io_output),
    .io_passthrough(mac_28_1_io_passthrough)
  );
  MAC mac_28_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_2_clock),
    .reset(mac_28_2_reset),
    .io_load(mac_28_2_io_load),
    .io_mulInput(mac_28_2_io_mulInput),
    .io_addInput(mac_28_2_io_addInput),
    .io_output(mac_28_2_io_output),
    .io_passthrough(mac_28_2_io_passthrough)
  );
  MAC mac_28_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_3_clock),
    .reset(mac_28_3_reset),
    .io_load(mac_28_3_io_load),
    .io_mulInput(mac_28_3_io_mulInput),
    .io_addInput(mac_28_3_io_addInput),
    .io_output(mac_28_3_io_output),
    .io_passthrough(mac_28_3_io_passthrough)
  );
  MAC mac_28_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_4_clock),
    .reset(mac_28_4_reset),
    .io_load(mac_28_4_io_load),
    .io_mulInput(mac_28_4_io_mulInput),
    .io_addInput(mac_28_4_io_addInput),
    .io_output(mac_28_4_io_output),
    .io_passthrough(mac_28_4_io_passthrough)
  );
  MAC mac_28_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_5_clock),
    .reset(mac_28_5_reset),
    .io_load(mac_28_5_io_load),
    .io_mulInput(mac_28_5_io_mulInput),
    .io_addInput(mac_28_5_io_addInput),
    .io_output(mac_28_5_io_output),
    .io_passthrough(mac_28_5_io_passthrough)
  );
  MAC mac_28_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_6_clock),
    .reset(mac_28_6_reset),
    .io_load(mac_28_6_io_load),
    .io_mulInput(mac_28_6_io_mulInput),
    .io_addInput(mac_28_6_io_addInput),
    .io_output(mac_28_6_io_output),
    .io_passthrough(mac_28_6_io_passthrough)
  );
  MAC mac_28_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_7_clock),
    .reset(mac_28_7_reset),
    .io_load(mac_28_7_io_load),
    .io_mulInput(mac_28_7_io_mulInput),
    .io_addInput(mac_28_7_io_addInput),
    .io_output(mac_28_7_io_output),
    .io_passthrough(mac_28_7_io_passthrough)
  );
  MAC mac_28_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_8_clock),
    .reset(mac_28_8_reset),
    .io_load(mac_28_8_io_load),
    .io_mulInput(mac_28_8_io_mulInput),
    .io_addInput(mac_28_8_io_addInput),
    .io_output(mac_28_8_io_output),
    .io_passthrough(mac_28_8_io_passthrough)
  );
  MAC mac_28_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_9_clock),
    .reset(mac_28_9_reset),
    .io_load(mac_28_9_io_load),
    .io_mulInput(mac_28_9_io_mulInput),
    .io_addInput(mac_28_9_io_addInput),
    .io_output(mac_28_9_io_output),
    .io_passthrough(mac_28_9_io_passthrough)
  );
  MAC mac_28_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_10_clock),
    .reset(mac_28_10_reset),
    .io_load(mac_28_10_io_load),
    .io_mulInput(mac_28_10_io_mulInput),
    .io_addInput(mac_28_10_io_addInput),
    .io_output(mac_28_10_io_output),
    .io_passthrough(mac_28_10_io_passthrough)
  );
  MAC mac_28_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_11_clock),
    .reset(mac_28_11_reset),
    .io_load(mac_28_11_io_load),
    .io_mulInput(mac_28_11_io_mulInput),
    .io_addInput(mac_28_11_io_addInput),
    .io_output(mac_28_11_io_output),
    .io_passthrough(mac_28_11_io_passthrough)
  );
  MAC mac_28_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_12_clock),
    .reset(mac_28_12_reset),
    .io_load(mac_28_12_io_load),
    .io_mulInput(mac_28_12_io_mulInput),
    .io_addInput(mac_28_12_io_addInput),
    .io_output(mac_28_12_io_output),
    .io_passthrough(mac_28_12_io_passthrough)
  );
  MAC mac_28_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_13_clock),
    .reset(mac_28_13_reset),
    .io_load(mac_28_13_io_load),
    .io_mulInput(mac_28_13_io_mulInput),
    .io_addInput(mac_28_13_io_addInput),
    .io_output(mac_28_13_io_output),
    .io_passthrough(mac_28_13_io_passthrough)
  );
  MAC mac_28_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_14_clock),
    .reset(mac_28_14_reset),
    .io_load(mac_28_14_io_load),
    .io_mulInput(mac_28_14_io_mulInput),
    .io_addInput(mac_28_14_io_addInput),
    .io_output(mac_28_14_io_output),
    .io_passthrough(mac_28_14_io_passthrough)
  );
  MAC mac_28_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_15_clock),
    .reset(mac_28_15_reset),
    .io_load(mac_28_15_io_load),
    .io_mulInput(mac_28_15_io_mulInput),
    .io_addInput(mac_28_15_io_addInput),
    .io_output(mac_28_15_io_output),
    .io_passthrough(mac_28_15_io_passthrough)
  );
  MAC mac_28_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_16_clock),
    .reset(mac_28_16_reset),
    .io_load(mac_28_16_io_load),
    .io_mulInput(mac_28_16_io_mulInput),
    .io_addInput(mac_28_16_io_addInput),
    .io_output(mac_28_16_io_output),
    .io_passthrough(mac_28_16_io_passthrough)
  );
  MAC mac_28_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_17_clock),
    .reset(mac_28_17_reset),
    .io_load(mac_28_17_io_load),
    .io_mulInput(mac_28_17_io_mulInput),
    .io_addInput(mac_28_17_io_addInput),
    .io_output(mac_28_17_io_output),
    .io_passthrough(mac_28_17_io_passthrough)
  );
  MAC mac_28_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_18_clock),
    .reset(mac_28_18_reset),
    .io_load(mac_28_18_io_load),
    .io_mulInput(mac_28_18_io_mulInput),
    .io_addInput(mac_28_18_io_addInput),
    .io_output(mac_28_18_io_output),
    .io_passthrough(mac_28_18_io_passthrough)
  );
  MAC mac_28_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_19_clock),
    .reset(mac_28_19_reset),
    .io_load(mac_28_19_io_load),
    .io_mulInput(mac_28_19_io_mulInput),
    .io_addInput(mac_28_19_io_addInput),
    .io_output(mac_28_19_io_output),
    .io_passthrough(mac_28_19_io_passthrough)
  );
  MAC mac_28_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_20_clock),
    .reset(mac_28_20_reset),
    .io_load(mac_28_20_io_load),
    .io_mulInput(mac_28_20_io_mulInput),
    .io_addInput(mac_28_20_io_addInput),
    .io_output(mac_28_20_io_output),
    .io_passthrough(mac_28_20_io_passthrough)
  );
  MAC mac_28_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_21_clock),
    .reset(mac_28_21_reset),
    .io_load(mac_28_21_io_load),
    .io_mulInput(mac_28_21_io_mulInput),
    .io_addInput(mac_28_21_io_addInput),
    .io_output(mac_28_21_io_output),
    .io_passthrough(mac_28_21_io_passthrough)
  );
  MAC mac_28_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_22_clock),
    .reset(mac_28_22_reset),
    .io_load(mac_28_22_io_load),
    .io_mulInput(mac_28_22_io_mulInput),
    .io_addInput(mac_28_22_io_addInput),
    .io_output(mac_28_22_io_output),
    .io_passthrough(mac_28_22_io_passthrough)
  );
  MAC mac_28_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_23_clock),
    .reset(mac_28_23_reset),
    .io_load(mac_28_23_io_load),
    .io_mulInput(mac_28_23_io_mulInput),
    .io_addInput(mac_28_23_io_addInput),
    .io_output(mac_28_23_io_output),
    .io_passthrough(mac_28_23_io_passthrough)
  );
  MAC mac_28_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_24_clock),
    .reset(mac_28_24_reset),
    .io_load(mac_28_24_io_load),
    .io_mulInput(mac_28_24_io_mulInput),
    .io_addInput(mac_28_24_io_addInput),
    .io_output(mac_28_24_io_output),
    .io_passthrough(mac_28_24_io_passthrough)
  );
  MAC mac_28_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_25_clock),
    .reset(mac_28_25_reset),
    .io_load(mac_28_25_io_load),
    .io_mulInput(mac_28_25_io_mulInput),
    .io_addInput(mac_28_25_io_addInput),
    .io_output(mac_28_25_io_output),
    .io_passthrough(mac_28_25_io_passthrough)
  );
  MAC mac_28_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_26_clock),
    .reset(mac_28_26_reset),
    .io_load(mac_28_26_io_load),
    .io_mulInput(mac_28_26_io_mulInput),
    .io_addInput(mac_28_26_io_addInput),
    .io_output(mac_28_26_io_output),
    .io_passthrough(mac_28_26_io_passthrough)
  );
  MAC mac_28_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_27_clock),
    .reset(mac_28_27_reset),
    .io_load(mac_28_27_io_load),
    .io_mulInput(mac_28_27_io_mulInput),
    .io_addInput(mac_28_27_io_addInput),
    .io_output(mac_28_27_io_output),
    .io_passthrough(mac_28_27_io_passthrough)
  );
  MAC mac_28_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_28_clock),
    .reset(mac_28_28_reset),
    .io_load(mac_28_28_io_load),
    .io_mulInput(mac_28_28_io_mulInput),
    .io_addInput(mac_28_28_io_addInput),
    .io_output(mac_28_28_io_output),
    .io_passthrough(mac_28_28_io_passthrough)
  );
  MAC mac_28_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_29_clock),
    .reset(mac_28_29_reset),
    .io_load(mac_28_29_io_load),
    .io_mulInput(mac_28_29_io_mulInput),
    .io_addInput(mac_28_29_io_addInput),
    .io_output(mac_28_29_io_output),
    .io_passthrough(mac_28_29_io_passthrough)
  );
  MAC mac_28_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_30_clock),
    .reset(mac_28_30_reset),
    .io_load(mac_28_30_io_load),
    .io_mulInput(mac_28_30_io_mulInput),
    .io_addInput(mac_28_30_io_addInput),
    .io_output(mac_28_30_io_output),
    .io_passthrough(mac_28_30_io_passthrough)
  );
  MAC mac_28_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_28_31_clock),
    .reset(mac_28_31_reset),
    .io_load(mac_28_31_io_load),
    .io_mulInput(mac_28_31_io_mulInput),
    .io_addInput(mac_28_31_io_addInput),
    .io_output(mac_28_31_io_output),
    .io_passthrough(mac_28_31_io_passthrough)
  );
  MAC mac_29_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_0_clock),
    .reset(mac_29_0_reset),
    .io_load(mac_29_0_io_load),
    .io_mulInput(mac_29_0_io_mulInput),
    .io_addInput(mac_29_0_io_addInput),
    .io_output(mac_29_0_io_output),
    .io_passthrough(mac_29_0_io_passthrough)
  );
  MAC mac_29_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_1_clock),
    .reset(mac_29_1_reset),
    .io_load(mac_29_1_io_load),
    .io_mulInput(mac_29_1_io_mulInput),
    .io_addInput(mac_29_1_io_addInput),
    .io_output(mac_29_1_io_output),
    .io_passthrough(mac_29_1_io_passthrough)
  );
  MAC mac_29_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_2_clock),
    .reset(mac_29_2_reset),
    .io_load(mac_29_2_io_load),
    .io_mulInput(mac_29_2_io_mulInput),
    .io_addInput(mac_29_2_io_addInput),
    .io_output(mac_29_2_io_output),
    .io_passthrough(mac_29_2_io_passthrough)
  );
  MAC mac_29_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_3_clock),
    .reset(mac_29_3_reset),
    .io_load(mac_29_3_io_load),
    .io_mulInput(mac_29_3_io_mulInput),
    .io_addInput(mac_29_3_io_addInput),
    .io_output(mac_29_3_io_output),
    .io_passthrough(mac_29_3_io_passthrough)
  );
  MAC mac_29_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_4_clock),
    .reset(mac_29_4_reset),
    .io_load(mac_29_4_io_load),
    .io_mulInput(mac_29_4_io_mulInput),
    .io_addInput(mac_29_4_io_addInput),
    .io_output(mac_29_4_io_output),
    .io_passthrough(mac_29_4_io_passthrough)
  );
  MAC mac_29_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_5_clock),
    .reset(mac_29_5_reset),
    .io_load(mac_29_5_io_load),
    .io_mulInput(mac_29_5_io_mulInput),
    .io_addInput(mac_29_5_io_addInput),
    .io_output(mac_29_5_io_output),
    .io_passthrough(mac_29_5_io_passthrough)
  );
  MAC mac_29_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_6_clock),
    .reset(mac_29_6_reset),
    .io_load(mac_29_6_io_load),
    .io_mulInput(mac_29_6_io_mulInput),
    .io_addInput(mac_29_6_io_addInput),
    .io_output(mac_29_6_io_output),
    .io_passthrough(mac_29_6_io_passthrough)
  );
  MAC mac_29_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_7_clock),
    .reset(mac_29_7_reset),
    .io_load(mac_29_7_io_load),
    .io_mulInput(mac_29_7_io_mulInput),
    .io_addInput(mac_29_7_io_addInput),
    .io_output(mac_29_7_io_output),
    .io_passthrough(mac_29_7_io_passthrough)
  );
  MAC mac_29_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_8_clock),
    .reset(mac_29_8_reset),
    .io_load(mac_29_8_io_load),
    .io_mulInput(mac_29_8_io_mulInput),
    .io_addInput(mac_29_8_io_addInput),
    .io_output(mac_29_8_io_output),
    .io_passthrough(mac_29_8_io_passthrough)
  );
  MAC mac_29_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_9_clock),
    .reset(mac_29_9_reset),
    .io_load(mac_29_9_io_load),
    .io_mulInput(mac_29_9_io_mulInput),
    .io_addInput(mac_29_9_io_addInput),
    .io_output(mac_29_9_io_output),
    .io_passthrough(mac_29_9_io_passthrough)
  );
  MAC mac_29_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_10_clock),
    .reset(mac_29_10_reset),
    .io_load(mac_29_10_io_load),
    .io_mulInput(mac_29_10_io_mulInput),
    .io_addInput(mac_29_10_io_addInput),
    .io_output(mac_29_10_io_output),
    .io_passthrough(mac_29_10_io_passthrough)
  );
  MAC mac_29_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_11_clock),
    .reset(mac_29_11_reset),
    .io_load(mac_29_11_io_load),
    .io_mulInput(mac_29_11_io_mulInput),
    .io_addInput(mac_29_11_io_addInput),
    .io_output(mac_29_11_io_output),
    .io_passthrough(mac_29_11_io_passthrough)
  );
  MAC mac_29_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_12_clock),
    .reset(mac_29_12_reset),
    .io_load(mac_29_12_io_load),
    .io_mulInput(mac_29_12_io_mulInput),
    .io_addInput(mac_29_12_io_addInput),
    .io_output(mac_29_12_io_output),
    .io_passthrough(mac_29_12_io_passthrough)
  );
  MAC mac_29_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_13_clock),
    .reset(mac_29_13_reset),
    .io_load(mac_29_13_io_load),
    .io_mulInput(mac_29_13_io_mulInput),
    .io_addInput(mac_29_13_io_addInput),
    .io_output(mac_29_13_io_output),
    .io_passthrough(mac_29_13_io_passthrough)
  );
  MAC mac_29_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_14_clock),
    .reset(mac_29_14_reset),
    .io_load(mac_29_14_io_load),
    .io_mulInput(mac_29_14_io_mulInput),
    .io_addInput(mac_29_14_io_addInput),
    .io_output(mac_29_14_io_output),
    .io_passthrough(mac_29_14_io_passthrough)
  );
  MAC mac_29_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_15_clock),
    .reset(mac_29_15_reset),
    .io_load(mac_29_15_io_load),
    .io_mulInput(mac_29_15_io_mulInput),
    .io_addInput(mac_29_15_io_addInput),
    .io_output(mac_29_15_io_output),
    .io_passthrough(mac_29_15_io_passthrough)
  );
  MAC mac_29_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_16_clock),
    .reset(mac_29_16_reset),
    .io_load(mac_29_16_io_load),
    .io_mulInput(mac_29_16_io_mulInput),
    .io_addInput(mac_29_16_io_addInput),
    .io_output(mac_29_16_io_output),
    .io_passthrough(mac_29_16_io_passthrough)
  );
  MAC mac_29_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_17_clock),
    .reset(mac_29_17_reset),
    .io_load(mac_29_17_io_load),
    .io_mulInput(mac_29_17_io_mulInput),
    .io_addInput(mac_29_17_io_addInput),
    .io_output(mac_29_17_io_output),
    .io_passthrough(mac_29_17_io_passthrough)
  );
  MAC mac_29_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_18_clock),
    .reset(mac_29_18_reset),
    .io_load(mac_29_18_io_load),
    .io_mulInput(mac_29_18_io_mulInput),
    .io_addInput(mac_29_18_io_addInput),
    .io_output(mac_29_18_io_output),
    .io_passthrough(mac_29_18_io_passthrough)
  );
  MAC mac_29_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_19_clock),
    .reset(mac_29_19_reset),
    .io_load(mac_29_19_io_load),
    .io_mulInput(mac_29_19_io_mulInput),
    .io_addInput(mac_29_19_io_addInput),
    .io_output(mac_29_19_io_output),
    .io_passthrough(mac_29_19_io_passthrough)
  );
  MAC mac_29_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_20_clock),
    .reset(mac_29_20_reset),
    .io_load(mac_29_20_io_load),
    .io_mulInput(mac_29_20_io_mulInput),
    .io_addInput(mac_29_20_io_addInput),
    .io_output(mac_29_20_io_output),
    .io_passthrough(mac_29_20_io_passthrough)
  );
  MAC mac_29_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_21_clock),
    .reset(mac_29_21_reset),
    .io_load(mac_29_21_io_load),
    .io_mulInput(mac_29_21_io_mulInput),
    .io_addInput(mac_29_21_io_addInput),
    .io_output(mac_29_21_io_output),
    .io_passthrough(mac_29_21_io_passthrough)
  );
  MAC mac_29_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_22_clock),
    .reset(mac_29_22_reset),
    .io_load(mac_29_22_io_load),
    .io_mulInput(mac_29_22_io_mulInput),
    .io_addInput(mac_29_22_io_addInput),
    .io_output(mac_29_22_io_output),
    .io_passthrough(mac_29_22_io_passthrough)
  );
  MAC mac_29_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_23_clock),
    .reset(mac_29_23_reset),
    .io_load(mac_29_23_io_load),
    .io_mulInput(mac_29_23_io_mulInput),
    .io_addInput(mac_29_23_io_addInput),
    .io_output(mac_29_23_io_output),
    .io_passthrough(mac_29_23_io_passthrough)
  );
  MAC mac_29_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_24_clock),
    .reset(mac_29_24_reset),
    .io_load(mac_29_24_io_load),
    .io_mulInput(mac_29_24_io_mulInput),
    .io_addInput(mac_29_24_io_addInput),
    .io_output(mac_29_24_io_output),
    .io_passthrough(mac_29_24_io_passthrough)
  );
  MAC mac_29_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_25_clock),
    .reset(mac_29_25_reset),
    .io_load(mac_29_25_io_load),
    .io_mulInput(mac_29_25_io_mulInput),
    .io_addInput(mac_29_25_io_addInput),
    .io_output(mac_29_25_io_output),
    .io_passthrough(mac_29_25_io_passthrough)
  );
  MAC mac_29_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_26_clock),
    .reset(mac_29_26_reset),
    .io_load(mac_29_26_io_load),
    .io_mulInput(mac_29_26_io_mulInput),
    .io_addInput(mac_29_26_io_addInput),
    .io_output(mac_29_26_io_output),
    .io_passthrough(mac_29_26_io_passthrough)
  );
  MAC mac_29_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_27_clock),
    .reset(mac_29_27_reset),
    .io_load(mac_29_27_io_load),
    .io_mulInput(mac_29_27_io_mulInput),
    .io_addInput(mac_29_27_io_addInput),
    .io_output(mac_29_27_io_output),
    .io_passthrough(mac_29_27_io_passthrough)
  );
  MAC mac_29_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_28_clock),
    .reset(mac_29_28_reset),
    .io_load(mac_29_28_io_load),
    .io_mulInput(mac_29_28_io_mulInput),
    .io_addInput(mac_29_28_io_addInput),
    .io_output(mac_29_28_io_output),
    .io_passthrough(mac_29_28_io_passthrough)
  );
  MAC mac_29_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_29_clock),
    .reset(mac_29_29_reset),
    .io_load(mac_29_29_io_load),
    .io_mulInput(mac_29_29_io_mulInput),
    .io_addInput(mac_29_29_io_addInput),
    .io_output(mac_29_29_io_output),
    .io_passthrough(mac_29_29_io_passthrough)
  );
  MAC mac_29_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_30_clock),
    .reset(mac_29_30_reset),
    .io_load(mac_29_30_io_load),
    .io_mulInput(mac_29_30_io_mulInput),
    .io_addInput(mac_29_30_io_addInput),
    .io_output(mac_29_30_io_output),
    .io_passthrough(mac_29_30_io_passthrough)
  );
  MAC mac_29_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_29_31_clock),
    .reset(mac_29_31_reset),
    .io_load(mac_29_31_io_load),
    .io_mulInput(mac_29_31_io_mulInput),
    .io_addInput(mac_29_31_io_addInput),
    .io_output(mac_29_31_io_output),
    .io_passthrough(mac_29_31_io_passthrough)
  );
  MAC mac_30_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_0_clock),
    .reset(mac_30_0_reset),
    .io_load(mac_30_0_io_load),
    .io_mulInput(mac_30_0_io_mulInput),
    .io_addInput(mac_30_0_io_addInput),
    .io_output(mac_30_0_io_output),
    .io_passthrough(mac_30_0_io_passthrough)
  );
  MAC mac_30_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_1_clock),
    .reset(mac_30_1_reset),
    .io_load(mac_30_1_io_load),
    .io_mulInput(mac_30_1_io_mulInput),
    .io_addInput(mac_30_1_io_addInput),
    .io_output(mac_30_1_io_output),
    .io_passthrough(mac_30_1_io_passthrough)
  );
  MAC mac_30_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_2_clock),
    .reset(mac_30_2_reset),
    .io_load(mac_30_2_io_load),
    .io_mulInput(mac_30_2_io_mulInput),
    .io_addInput(mac_30_2_io_addInput),
    .io_output(mac_30_2_io_output),
    .io_passthrough(mac_30_2_io_passthrough)
  );
  MAC mac_30_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_3_clock),
    .reset(mac_30_3_reset),
    .io_load(mac_30_3_io_load),
    .io_mulInput(mac_30_3_io_mulInput),
    .io_addInput(mac_30_3_io_addInput),
    .io_output(mac_30_3_io_output),
    .io_passthrough(mac_30_3_io_passthrough)
  );
  MAC mac_30_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_4_clock),
    .reset(mac_30_4_reset),
    .io_load(mac_30_4_io_load),
    .io_mulInput(mac_30_4_io_mulInput),
    .io_addInput(mac_30_4_io_addInput),
    .io_output(mac_30_4_io_output),
    .io_passthrough(mac_30_4_io_passthrough)
  );
  MAC mac_30_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_5_clock),
    .reset(mac_30_5_reset),
    .io_load(mac_30_5_io_load),
    .io_mulInput(mac_30_5_io_mulInput),
    .io_addInput(mac_30_5_io_addInput),
    .io_output(mac_30_5_io_output),
    .io_passthrough(mac_30_5_io_passthrough)
  );
  MAC mac_30_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_6_clock),
    .reset(mac_30_6_reset),
    .io_load(mac_30_6_io_load),
    .io_mulInput(mac_30_6_io_mulInput),
    .io_addInput(mac_30_6_io_addInput),
    .io_output(mac_30_6_io_output),
    .io_passthrough(mac_30_6_io_passthrough)
  );
  MAC mac_30_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_7_clock),
    .reset(mac_30_7_reset),
    .io_load(mac_30_7_io_load),
    .io_mulInput(mac_30_7_io_mulInput),
    .io_addInput(mac_30_7_io_addInput),
    .io_output(mac_30_7_io_output),
    .io_passthrough(mac_30_7_io_passthrough)
  );
  MAC mac_30_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_8_clock),
    .reset(mac_30_8_reset),
    .io_load(mac_30_8_io_load),
    .io_mulInput(mac_30_8_io_mulInput),
    .io_addInput(mac_30_8_io_addInput),
    .io_output(mac_30_8_io_output),
    .io_passthrough(mac_30_8_io_passthrough)
  );
  MAC mac_30_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_9_clock),
    .reset(mac_30_9_reset),
    .io_load(mac_30_9_io_load),
    .io_mulInput(mac_30_9_io_mulInput),
    .io_addInput(mac_30_9_io_addInput),
    .io_output(mac_30_9_io_output),
    .io_passthrough(mac_30_9_io_passthrough)
  );
  MAC mac_30_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_10_clock),
    .reset(mac_30_10_reset),
    .io_load(mac_30_10_io_load),
    .io_mulInput(mac_30_10_io_mulInput),
    .io_addInput(mac_30_10_io_addInput),
    .io_output(mac_30_10_io_output),
    .io_passthrough(mac_30_10_io_passthrough)
  );
  MAC mac_30_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_11_clock),
    .reset(mac_30_11_reset),
    .io_load(mac_30_11_io_load),
    .io_mulInput(mac_30_11_io_mulInput),
    .io_addInput(mac_30_11_io_addInput),
    .io_output(mac_30_11_io_output),
    .io_passthrough(mac_30_11_io_passthrough)
  );
  MAC mac_30_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_12_clock),
    .reset(mac_30_12_reset),
    .io_load(mac_30_12_io_load),
    .io_mulInput(mac_30_12_io_mulInput),
    .io_addInput(mac_30_12_io_addInput),
    .io_output(mac_30_12_io_output),
    .io_passthrough(mac_30_12_io_passthrough)
  );
  MAC mac_30_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_13_clock),
    .reset(mac_30_13_reset),
    .io_load(mac_30_13_io_load),
    .io_mulInput(mac_30_13_io_mulInput),
    .io_addInput(mac_30_13_io_addInput),
    .io_output(mac_30_13_io_output),
    .io_passthrough(mac_30_13_io_passthrough)
  );
  MAC mac_30_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_14_clock),
    .reset(mac_30_14_reset),
    .io_load(mac_30_14_io_load),
    .io_mulInput(mac_30_14_io_mulInput),
    .io_addInput(mac_30_14_io_addInput),
    .io_output(mac_30_14_io_output),
    .io_passthrough(mac_30_14_io_passthrough)
  );
  MAC mac_30_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_15_clock),
    .reset(mac_30_15_reset),
    .io_load(mac_30_15_io_load),
    .io_mulInput(mac_30_15_io_mulInput),
    .io_addInput(mac_30_15_io_addInput),
    .io_output(mac_30_15_io_output),
    .io_passthrough(mac_30_15_io_passthrough)
  );
  MAC mac_30_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_16_clock),
    .reset(mac_30_16_reset),
    .io_load(mac_30_16_io_load),
    .io_mulInput(mac_30_16_io_mulInput),
    .io_addInput(mac_30_16_io_addInput),
    .io_output(mac_30_16_io_output),
    .io_passthrough(mac_30_16_io_passthrough)
  );
  MAC mac_30_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_17_clock),
    .reset(mac_30_17_reset),
    .io_load(mac_30_17_io_load),
    .io_mulInput(mac_30_17_io_mulInput),
    .io_addInput(mac_30_17_io_addInput),
    .io_output(mac_30_17_io_output),
    .io_passthrough(mac_30_17_io_passthrough)
  );
  MAC mac_30_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_18_clock),
    .reset(mac_30_18_reset),
    .io_load(mac_30_18_io_load),
    .io_mulInput(mac_30_18_io_mulInput),
    .io_addInput(mac_30_18_io_addInput),
    .io_output(mac_30_18_io_output),
    .io_passthrough(mac_30_18_io_passthrough)
  );
  MAC mac_30_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_19_clock),
    .reset(mac_30_19_reset),
    .io_load(mac_30_19_io_load),
    .io_mulInput(mac_30_19_io_mulInput),
    .io_addInput(mac_30_19_io_addInput),
    .io_output(mac_30_19_io_output),
    .io_passthrough(mac_30_19_io_passthrough)
  );
  MAC mac_30_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_20_clock),
    .reset(mac_30_20_reset),
    .io_load(mac_30_20_io_load),
    .io_mulInput(mac_30_20_io_mulInput),
    .io_addInput(mac_30_20_io_addInput),
    .io_output(mac_30_20_io_output),
    .io_passthrough(mac_30_20_io_passthrough)
  );
  MAC mac_30_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_21_clock),
    .reset(mac_30_21_reset),
    .io_load(mac_30_21_io_load),
    .io_mulInput(mac_30_21_io_mulInput),
    .io_addInput(mac_30_21_io_addInput),
    .io_output(mac_30_21_io_output),
    .io_passthrough(mac_30_21_io_passthrough)
  );
  MAC mac_30_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_22_clock),
    .reset(mac_30_22_reset),
    .io_load(mac_30_22_io_load),
    .io_mulInput(mac_30_22_io_mulInput),
    .io_addInput(mac_30_22_io_addInput),
    .io_output(mac_30_22_io_output),
    .io_passthrough(mac_30_22_io_passthrough)
  );
  MAC mac_30_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_23_clock),
    .reset(mac_30_23_reset),
    .io_load(mac_30_23_io_load),
    .io_mulInput(mac_30_23_io_mulInput),
    .io_addInput(mac_30_23_io_addInput),
    .io_output(mac_30_23_io_output),
    .io_passthrough(mac_30_23_io_passthrough)
  );
  MAC mac_30_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_24_clock),
    .reset(mac_30_24_reset),
    .io_load(mac_30_24_io_load),
    .io_mulInput(mac_30_24_io_mulInput),
    .io_addInput(mac_30_24_io_addInput),
    .io_output(mac_30_24_io_output),
    .io_passthrough(mac_30_24_io_passthrough)
  );
  MAC mac_30_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_25_clock),
    .reset(mac_30_25_reset),
    .io_load(mac_30_25_io_load),
    .io_mulInput(mac_30_25_io_mulInput),
    .io_addInput(mac_30_25_io_addInput),
    .io_output(mac_30_25_io_output),
    .io_passthrough(mac_30_25_io_passthrough)
  );
  MAC mac_30_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_26_clock),
    .reset(mac_30_26_reset),
    .io_load(mac_30_26_io_load),
    .io_mulInput(mac_30_26_io_mulInput),
    .io_addInput(mac_30_26_io_addInput),
    .io_output(mac_30_26_io_output),
    .io_passthrough(mac_30_26_io_passthrough)
  );
  MAC mac_30_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_27_clock),
    .reset(mac_30_27_reset),
    .io_load(mac_30_27_io_load),
    .io_mulInput(mac_30_27_io_mulInput),
    .io_addInput(mac_30_27_io_addInput),
    .io_output(mac_30_27_io_output),
    .io_passthrough(mac_30_27_io_passthrough)
  );
  MAC mac_30_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_28_clock),
    .reset(mac_30_28_reset),
    .io_load(mac_30_28_io_load),
    .io_mulInput(mac_30_28_io_mulInput),
    .io_addInput(mac_30_28_io_addInput),
    .io_output(mac_30_28_io_output),
    .io_passthrough(mac_30_28_io_passthrough)
  );
  MAC mac_30_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_29_clock),
    .reset(mac_30_29_reset),
    .io_load(mac_30_29_io_load),
    .io_mulInput(mac_30_29_io_mulInput),
    .io_addInput(mac_30_29_io_addInput),
    .io_output(mac_30_29_io_output),
    .io_passthrough(mac_30_29_io_passthrough)
  );
  MAC mac_30_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_30_clock),
    .reset(mac_30_30_reset),
    .io_load(mac_30_30_io_load),
    .io_mulInput(mac_30_30_io_mulInput),
    .io_addInput(mac_30_30_io_addInput),
    .io_output(mac_30_30_io_output),
    .io_passthrough(mac_30_30_io_passthrough)
  );
  MAC mac_30_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_30_31_clock),
    .reset(mac_30_31_reset),
    .io_load(mac_30_31_io_load),
    .io_mulInput(mac_30_31_io_mulInput),
    .io_addInput(mac_30_31_io_addInput),
    .io_output(mac_30_31_io_output),
    .io_passthrough(mac_30_31_io_passthrough)
  );
  MAC mac_31_0 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_0_clock),
    .reset(mac_31_0_reset),
    .io_load(mac_31_0_io_load),
    .io_mulInput(mac_31_0_io_mulInput),
    .io_addInput(mac_31_0_io_addInput),
    .io_output(mac_31_0_io_output),
    .io_passthrough(mac_31_0_io_passthrough)
  );
  MAC mac_31_1 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_1_clock),
    .reset(mac_31_1_reset),
    .io_load(mac_31_1_io_load),
    .io_mulInput(mac_31_1_io_mulInput),
    .io_addInput(mac_31_1_io_addInput),
    .io_output(mac_31_1_io_output),
    .io_passthrough(mac_31_1_io_passthrough)
  );
  MAC mac_31_2 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_2_clock),
    .reset(mac_31_2_reset),
    .io_load(mac_31_2_io_load),
    .io_mulInput(mac_31_2_io_mulInput),
    .io_addInput(mac_31_2_io_addInput),
    .io_output(mac_31_2_io_output),
    .io_passthrough(mac_31_2_io_passthrough)
  );
  MAC mac_31_3 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_3_clock),
    .reset(mac_31_3_reset),
    .io_load(mac_31_3_io_load),
    .io_mulInput(mac_31_3_io_mulInput),
    .io_addInput(mac_31_3_io_addInput),
    .io_output(mac_31_3_io_output),
    .io_passthrough(mac_31_3_io_passthrough)
  );
  MAC mac_31_4 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_4_clock),
    .reset(mac_31_4_reset),
    .io_load(mac_31_4_io_load),
    .io_mulInput(mac_31_4_io_mulInput),
    .io_addInput(mac_31_4_io_addInput),
    .io_output(mac_31_4_io_output),
    .io_passthrough(mac_31_4_io_passthrough)
  );
  MAC mac_31_5 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_5_clock),
    .reset(mac_31_5_reset),
    .io_load(mac_31_5_io_load),
    .io_mulInput(mac_31_5_io_mulInput),
    .io_addInput(mac_31_5_io_addInput),
    .io_output(mac_31_5_io_output),
    .io_passthrough(mac_31_5_io_passthrough)
  );
  MAC mac_31_6 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_6_clock),
    .reset(mac_31_6_reset),
    .io_load(mac_31_6_io_load),
    .io_mulInput(mac_31_6_io_mulInput),
    .io_addInput(mac_31_6_io_addInput),
    .io_output(mac_31_6_io_output),
    .io_passthrough(mac_31_6_io_passthrough)
  );
  MAC mac_31_7 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_7_clock),
    .reset(mac_31_7_reset),
    .io_load(mac_31_7_io_load),
    .io_mulInput(mac_31_7_io_mulInput),
    .io_addInput(mac_31_7_io_addInput),
    .io_output(mac_31_7_io_output),
    .io_passthrough(mac_31_7_io_passthrough)
  );
  MAC mac_31_8 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_8_clock),
    .reset(mac_31_8_reset),
    .io_load(mac_31_8_io_load),
    .io_mulInput(mac_31_8_io_mulInput),
    .io_addInput(mac_31_8_io_addInput),
    .io_output(mac_31_8_io_output),
    .io_passthrough(mac_31_8_io_passthrough)
  );
  MAC mac_31_9 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_9_clock),
    .reset(mac_31_9_reset),
    .io_load(mac_31_9_io_load),
    .io_mulInput(mac_31_9_io_mulInput),
    .io_addInput(mac_31_9_io_addInput),
    .io_output(mac_31_9_io_output),
    .io_passthrough(mac_31_9_io_passthrough)
  );
  MAC mac_31_10 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_10_clock),
    .reset(mac_31_10_reset),
    .io_load(mac_31_10_io_load),
    .io_mulInput(mac_31_10_io_mulInput),
    .io_addInput(mac_31_10_io_addInput),
    .io_output(mac_31_10_io_output),
    .io_passthrough(mac_31_10_io_passthrough)
  );
  MAC mac_31_11 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_11_clock),
    .reset(mac_31_11_reset),
    .io_load(mac_31_11_io_load),
    .io_mulInput(mac_31_11_io_mulInput),
    .io_addInput(mac_31_11_io_addInput),
    .io_output(mac_31_11_io_output),
    .io_passthrough(mac_31_11_io_passthrough)
  );
  MAC mac_31_12 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_12_clock),
    .reset(mac_31_12_reset),
    .io_load(mac_31_12_io_load),
    .io_mulInput(mac_31_12_io_mulInput),
    .io_addInput(mac_31_12_io_addInput),
    .io_output(mac_31_12_io_output),
    .io_passthrough(mac_31_12_io_passthrough)
  );
  MAC mac_31_13 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_13_clock),
    .reset(mac_31_13_reset),
    .io_load(mac_31_13_io_load),
    .io_mulInput(mac_31_13_io_mulInput),
    .io_addInput(mac_31_13_io_addInput),
    .io_output(mac_31_13_io_output),
    .io_passthrough(mac_31_13_io_passthrough)
  );
  MAC mac_31_14 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_14_clock),
    .reset(mac_31_14_reset),
    .io_load(mac_31_14_io_load),
    .io_mulInput(mac_31_14_io_mulInput),
    .io_addInput(mac_31_14_io_addInput),
    .io_output(mac_31_14_io_output),
    .io_passthrough(mac_31_14_io_passthrough)
  );
  MAC mac_31_15 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_15_clock),
    .reset(mac_31_15_reset),
    .io_load(mac_31_15_io_load),
    .io_mulInput(mac_31_15_io_mulInput),
    .io_addInput(mac_31_15_io_addInput),
    .io_output(mac_31_15_io_output),
    .io_passthrough(mac_31_15_io_passthrough)
  );
  MAC mac_31_16 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_16_clock),
    .reset(mac_31_16_reset),
    .io_load(mac_31_16_io_load),
    .io_mulInput(mac_31_16_io_mulInput),
    .io_addInput(mac_31_16_io_addInput),
    .io_output(mac_31_16_io_output),
    .io_passthrough(mac_31_16_io_passthrough)
  );
  MAC mac_31_17 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_17_clock),
    .reset(mac_31_17_reset),
    .io_load(mac_31_17_io_load),
    .io_mulInput(mac_31_17_io_mulInput),
    .io_addInput(mac_31_17_io_addInput),
    .io_output(mac_31_17_io_output),
    .io_passthrough(mac_31_17_io_passthrough)
  );
  MAC mac_31_18 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_18_clock),
    .reset(mac_31_18_reset),
    .io_load(mac_31_18_io_load),
    .io_mulInput(mac_31_18_io_mulInput),
    .io_addInput(mac_31_18_io_addInput),
    .io_output(mac_31_18_io_output),
    .io_passthrough(mac_31_18_io_passthrough)
  );
  MAC mac_31_19 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_19_clock),
    .reset(mac_31_19_reset),
    .io_load(mac_31_19_io_load),
    .io_mulInput(mac_31_19_io_mulInput),
    .io_addInput(mac_31_19_io_addInput),
    .io_output(mac_31_19_io_output),
    .io_passthrough(mac_31_19_io_passthrough)
  );
  MAC mac_31_20 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_20_clock),
    .reset(mac_31_20_reset),
    .io_load(mac_31_20_io_load),
    .io_mulInput(mac_31_20_io_mulInput),
    .io_addInput(mac_31_20_io_addInput),
    .io_output(mac_31_20_io_output),
    .io_passthrough(mac_31_20_io_passthrough)
  );
  MAC mac_31_21 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_21_clock),
    .reset(mac_31_21_reset),
    .io_load(mac_31_21_io_load),
    .io_mulInput(mac_31_21_io_mulInput),
    .io_addInput(mac_31_21_io_addInput),
    .io_output(mac_31_21_io_output),
    .io_passthrough(mac_31_21_io_passthrough)
  );
  MAC mac_31_22 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_22_clock),
    .reset(mac_31_22_reset),
    .io_load(mac_31_22_io_load),
    .io_mulInput(mac_31_22_io_mulInput),
    .io_addInput(mac_31_22_io_addInput),
    .io_output(mac_31_22_io_output),
    .io_passthrough(mac_31_22_io_passthrough)
  );
  MAC mac_31_23 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_23_clock),
    .reset(mac_31_23_reset),
    .io_load(mac_31_23_io_load),
    .io_mulInput(mac_31_23_io_mulInput),
    .io_addInput(mac_31_23_io_addInput),
    .io_output(mac_31_23_io_output),
    .io_passthrough(mac_31_23_io_passthrough)
  );
  MAC mac_31_24 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_24_clock),
    .reset(mac_31_24_reset),
    .io_load(mac_31_24_io_load),
    .io_mulInput(mac_31_24_io_mulInput),
    .io_addInput(mac_31_24_io_addInput),
    .io_output(mac_31_24_io_output),
    .io_passthrough(mac_31_24_io_passthrough)
  );
  MAC mac_31_25 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_25_clock),
    .reset(mac_31_25_reset),
    .io_load(mac_31_25_io_load),
    .io_mulInput(mac_31_25_io_mulInput),
    .io_addInput(mac_31_25_io_addInput),
    .io_output(mac_31_25_io_output),
    .io_passthrough(mac_31_25_io_passthrough)
  );
  MAC mac_31_26 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_26_clock),
    .reset(mac_31_26_reset),
    .io_load(mac_31_26_io_load),
    .io_mulInput(mac_31_26_io_mulInput),
    .io_addInput(mac_31_26_io_addInput),
    .io_output(mac_31_26_io_output),
    .io_passthrough(mac_31_26_io_passthrough)
  );
  MAC mac_31_27 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_27_clock),
    .reset(mac_31_27_reset),
    .io_load(mac_31_27_io_load),
    .io_mulInput(mac_31_27_io_mulInput),
    .io_addInput(mac_31_27_io_addInput),
    .io_output(mac_31_27_io_output),
    .io_passthrough(mac_31_27_io_passthrough)
  );
  MAC mac_31_28 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_28_clock),
    .reset(mac_31_28_reset),
    .io_load(mac_31_28_io_load),
    .io_mulInput(mac_31_28_io_mulInput),
    .io_addInput(mac_31_28_io_addInput),
    .io_output(mac_31_28_io_output),
    .io_passthrough(mac_31_28_io_passthrough)
  );
  MAC mac_31_29 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_29_clock),
    .reset(mac_31_29_reset),
    .io_load(mac_31_29_io_load),
    .io_mulInput(mac_31_29_io_mulInput),
    .io_addInput(mac_31_29_io_addInput),
    .io_output(mac_31_29_io_output),
    .io_passthrough(mac_31_29_io_passthrough)
  );
  MAC mac_31_30 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_30_clock),
    .reset(mac_31_30_reset),
    .io_load(mac_31_30_io_load),
    .io_mulInput(mac_31_30_io_mulInput),
    .io_addInput(mac_31_30_io_addInput),
    .io_output(mac_31_30_io_output),
    .io_passthrough(mac_31_30_io_passthrough)
  );
  MAC mac_31_31 ( // @[InnerSystolicArray.scala 34:50]
    .clock(mac_31_31_clock),
    .reset(mac_31_31_reset),
    .io_load(mac_31_31_io_load),
    .io_mulInput(mac_31_31_io_mulInput),
    .io_addInput(mac_31_31_io_addInput),
    .io_output(mac_31_31_io_output),
    .io_passthrough(mac_31_31_io_passthrough)
  );
  assign io_output_0 = io_output_0_sr_30; // @[InnerSystolicArray.scala 75:18]
  assign io_output_1 = io_output_1_sr_29; // @[InnerSystolicArray.scala 75:18]
  assign io_output_2 = io_output_2_sr_28; // @[InnerSystolicArray.scala 75:18]
  assign io_output_3 = io_output_3_sr_27; // @[InnerSystolicArray.scala 75:18]
  assign io_output_4 = io_output_4_sr_26; // @[InnerSystolicArray.scala 75:18]
  assign io_output_5 = io_output_5_sr_25; // @[InnerSystolicArray.scala 75:18]
  assign io_output_6 = io_output_6_sr_24; // @[InnerSystolicArray.scala 75:18]
  assign io_output_7 = io_output_7_sr_23; // @[InnerSystolicArray.scala 75:18]
  assign io_output_8 = io_output_8_sr_22; // @[InnerSystolicArray.scala 75:18]
  assign io_output_9 = io_output_9_sr_21; // @[InnerSystolicArray.scala 75:18]
  assign io_output_10 = io_output_10_sr_20; // @[InnerSystolicArray.scala 75:18]
  assign io_output_11 = io_output_11_sr_19; // @[InnerSystolicArray.scala 75:18]
  assign io_output_12 = io_output_12_sr_18; // @[InnerSystolicArray.scala 75:18]
  assign io_output_13 = io_output_13_sr_17; // @[InnerSystolicArray.scala 75:18]
  assign io_output_14 = io_output_14_sr_16; // @[InnerSystolicArray.scala 75:18]
  assign io_output_15 = io_output_15_sr_15; // @[InnerSystolicArray.scala 75:18]
  assign io_output_16 = io_output_16_sr_14; // @[InnerSystolicArray.scala 75:18]
  assign io_output_17 = io_output_17_sr_13; // @[InnerSystolicArray.scala 75:18]
  assign io_output_18 = io_output_18_sr_12; // @[InnerSystolicArray.scala 75:18]
  assign io_output_19 = io_output_19_sr_11; // @[InnerSystolicArray.scala 75:18]
  assign io_output_20 = io_output_20_sr_10; // @[InnerSystolicArray.scala 75:18]
  assign io_output_21 = io_output_21_sr_9; // @[InnerSystolicArray.scala 75:18]
  assign io_output_22 = io_output_22_sr_8; // @[InnerSystolicArray.scala 75:18]
  assign io_output_23 = io_output_23_sr_7; // @[InnerSystolicArray.scala 75:18]
  assign io_output_24 = io_output_24_sr_6; // @[InnerSystolicArray.scala 75:18]
  assign io_output_25 = io_output_25_sr_5; // @[InnerSystolicArray.scala 75:18]
  assign io_output_26 = io_output_26_sr_4; // @[InnerSystolicArray.scala 75:18]
  assign io_output_27 = io_output_27_sr_3; // @[InnerSystolicArray.scala 75:18]
  assign io_output_28 = io_output_28_sr_2; // @[InnerSystolicArray.scala 75:18]
  assign io_output_29 = io_output_29_sr_1; // @[InnerSystolicArray.scala 75:18]
  assign io_output_30 = io_output_30_sr_0; // @[InnerSystolicArray.scala 75:18]
  assign io_output_31 = mac_31_31_io_output; // @[InnerSystolicArray.scala 75:18]
  assign mac_0_0_clock = clock;
  assign mac_0_0_reset = reset;
  assign mac_0_0_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_0_io_mulInput = io_input_0; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_0_io_addInput = bias_0; // @[InnerSystolicArray.scala 57:27]
  assign mac_0_1_clock = clock;
  assign mac_0_1_reset = reset;
  assign mac_0_1_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_1_io_mulInput = mac_0_1_io_mulInput_sr_0; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_1_io_addInput = mac_0_0_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_2_clock = clock;
  assign mac_0_2_reset = reset;
  assign mac_0_2_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_2_io_mulInput = mac_0_2_io_mulInput_sr_1; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_2_io_addInput = mac_0_1_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_3_clock = clock;
  assign mac_0_3_reset = reset;
  assign mac_0_3_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_3_io_mulInput = mac_0_3_io_mulInput_sr_2; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_3_io_addInput = mac_0_2_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_4_clock = clock;
  assign mac_0_4_reset = reset;
  assign mac_0_4_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_4_io_mulInput = mac_0_4_io_mulInput_sr_3; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_4_io_addInput = mac_0_3_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_5_clock = clock;
  assign mac_0_5_reset = reset;
  assign mac_0_5_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_5_io_mulInput = mac_0_5_io_mulInput_sr_4; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_5_io_addInput = mac_0_4_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_6_clock = clock;
  assign mac_0_6_reset = reset;
  assign mac_0_6_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_6_io_mulInput = mac_0_6_io_mulInput_sr_5; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_6_io_addInput = mac_0_5_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_7_clock = clock;
  assign mac_0_7_reset = reset;
  assign mac_0_7_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_7_io_mulInput = mac_0_7_io_mulInput_sr_6; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_7_io_addInput = mac_0_6_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_8_clock = clock;
  assign mac_0_8_reset = reset;
  assign mac_0_8_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_8_io_mulInput = mac_0_8_io_mulInput_sr_7; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_8_io_addInput = mac_0_7_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_9_clock = clock;
  assign mac_0_9_reset = reset;
  assign mac_0_9_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_9_io_mulInput = mac_0_9_io_mulInput_sr_8; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_9_io_addInput = mac_0_8_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_10_clock = clock;
  assign mac_0_10_reset = reset;
  assign mac_0_10_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_10_io_mulInput = mac_0_10_io_mulInput_sr_9; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_10_io_addInput = mac_0_9_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_11_clock = clock;
  assign mac_0_11_reset = reset;
  assign mac_0_11_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_11_io_mulInput = mac_0_11_io_mulInput_sr_10; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_11_io_addInput = mac_0_10_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_12_clock = clock;
  assign mac_0_12_reset = reset;
  assign mac_0_12_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_12_io_mulInput = mac_0_12_io_mulInput_sr_11; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_12_io_addInput = mac_0_11_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_13_clock = clock;
  assign mac_0_13_reset = reset;
  assign mac_0_13_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_13_io_mulInput = mac_0_13_io_mulInput_sr_12; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_13_io_addInput = mac_0_12_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_14_clock = clock;
  assign mac_0_14_reset = reset;
  assign mac_0_14_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_14_io_mulInput = mac_0_14_io_mulInput_sr_13; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_14_io_addInput = mac_0_13_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_15_clock = clock;
  assign mac_0_15_reset = reset;
  assign mac_0_15_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_15_io_mulInput = mac_0_15_io_mulInput_sr_14; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_15_io_addInput = mac_0_14_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_16_clock = clock;
  assign mac_0_16_reset = reset;
  assign mac_0_16_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_16_io_mulInput = mac_0_16_io_mulInput_sr_15; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_16_io_addInput = mac_0_15_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_17_clock = clock;
  assign mac_0_17_reset = reset;
  assign mac_0_17_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_17_io_mulInput = mac_0_17_io_mulInput_sr_16; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_17_io_addInput = mac_0_16_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_18_clock = clock;
  assign mac_0_18_reset = reset;
  assign mac_0_18_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_18_io_mulInput = mac_0_18_io_mulInput_sr_17; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_18_io_addInput = mac_0_17_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_19_clock = clock;
  assign mac_0_19_reset = reset;
  assign mac_0_19_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_19_io_mulInput = mac_0_19_io_mulInput_sr_18; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_19_io_addInput = mac_0_18_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_20_clock = clock;
  assign mac_0_20_reset = reset;
  assign mac_0_20_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_20_io_mulInput = mac_0_20_io_mulInput_sr_19; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_20_io_addInput = mac_0_19_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_21_clock = clock;
  assign mac_0_21_reset = reset;
  assign mac_0_21_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_21_io_mulInput = mac_0_21_io_mulInput_sr_20; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_21_io_addInput = mac_0_20_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_22_clock = clock;
  assign mac_0_22_reset = reset;
  assign mac_0_22_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_22_io_mulInput = mac_0_22_io_mulInput_sr_21; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_22_io_addInput = mac_0_21_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_23_clock = clock;
  assign mac_0_23_reset = reset;
  assign mac_0_23_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_23_io_mulInput = mac_0_23_io_mulInput_sr_22; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_23_io_addInput = mac_0_22_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_24_clock = clock;
  assign mac_0_24_reset = reset;
  assign mac_0_24_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_24_io_mulInput = mac_0_24_io_mulInput_sr_23; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_24_io_addInput = mac_0_23_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_25_clock = clock;
  assign mac_0_25_reset = reset;
  assign mac_0_25_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_25_io_mulInput = mac_0_25_io_mulInput_sr_24; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_25_io_addInput = mac_0_24_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_26_clock = clock;
  assign mac_0_26_reset = reset;
  assign mac_0_26_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_26_io_mulInput = mac_0_26_io_mulInput_sr_25; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_26_io_addInput = mac_0_25_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_27_clock = clock;
  assign mac_0_27_reset = reset;
  assign mac_0_27_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_27_io_mulInput = mac_0_27_io_mulInput_sr_26; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_27_io_addInput = mac_0_26_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_28_clock = clock;
  assign mac_0_28_reset = reset;
  assign mac_0_28_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_28_io_mulInput = mac_0_28_io_mulInput_sr_27; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_28_io_addInput = mac_0_27_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_29_clock = clock;
  assign mac_0_29_reset = reset;
  assign mac_0_29_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_29_io_mulInput = mac_0_29_io_mulInput_sr_28; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_29_io_addInput = mac_0_28_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_30_clock = clock;
  assign mac_0_30_reset = reset;
  assign mac_0_30_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_30_io_mulInput = mac_0_30_io_mulInput_sr_29; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_30_io_addInput = mac_0_29_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_0_31_clock = clock;
  assign mac_0_31_reset = reset;
  assign mac_0_31_io_load = io_load; // @[InnerSystolicArray.scala 52:23]
  assign mac_0_31_io_mulInput = mac_0_31_io_mulInput_sr_30; // @[InnerSystolicArray.scala 48:27]
  assign mac_0_31_io_addInput = mac_0_30_io_output; // @[InnerSystolicArray.scala 50:29]
  assign mac_1_0_clock = clock;
  assign mac_1_0_reset = reset;
  assign mac_1_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_1_0_io_mulInput = mac_0_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_1_0_io_addInput = bias_1; // @[InnerSystolicArray.scala 57:27]
  assign mac_1_1_clock = clock;
  assign mac_1_1_reset = reset;
  assign mac_1_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_1_io_mulInput = mac_0_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_1_io_addInput = mac_1_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_2_clock = clock;
  assign mac_1_2_reset = reset;
  assign mac_1_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_2_io_mulInput = mac_0_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_2_io_addInput = mac_1_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_3_clock = clock;
  assign mac_1_3_reset = reset;
  assign mac_1_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_3_io_mulInput = mac_0_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_3_io_addInput = mac_1_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_4_clock = clock;
  assign mac_1_4_reset = reset;
  assign mac_1_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_4_io_mulInput = mac_0_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_4_io_addInput = mac_1_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_5_clock = clock;
  assign mac_1_5_reset = reset;
  assign mac_1_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_5_io_mulInput = mac_0_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_5_io_addInput = mac_1_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_6_clock = clock;
  assign mac_1_6_reset = reset;
  assign mac_1_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_6_io_mulInput = mac_0_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_6_io_addInput = mac_1_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_7_clock = clock;
  assign mac_1_7_reset = reset;
  assign mac_1_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_7_io_mulInput = mac_0_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_7_io_addInput = mac_1_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_8_clock = clock;
  assign mac_1_8_reset = reset;
  assign mac_1_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_8_io_mulInput = mac_0_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_8_io_addInput = mac_1_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_9_clock = clock;
  assign mac_1_9_reset = reset;
  assign mac_1_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_9_io_mulInput = mac_0_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_9_io_addInput = mac_1_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_10_clock = clock;
  assign mac_1_10_reset = reset;
  assign mac_1_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_10_io_mulInput = mac_0_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_10_io_addInput = mac_1_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_11_clock = clock;
  assign mac_1_11_reset = reset;
  assign mac_1_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_11_io_mulInput = mac_0_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_11_io_addInput = mac_1_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_12_clock = clock;
  assign mac_1_12_reset = reset;
  assign mac_1_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_12_io_mulInput = mac_0_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_12_io_addInput = mac_1_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_13_clock = clock;
  assign mac_1_13_reset = reset;
  assign mac_1_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_13_io_mulInput = mac_0_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_13_io_addInput = mac_1_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_14_clock = clock;
  assign mac_1_14_reset = reset;
  assign mac_1_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_14_io_mulInput = mac_0_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_14_io_addInput = mac_1_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_15_clock = clock;
  assign mac_1_15_reset = reset;
  assign mac_1_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_15_io_mulInput = mac_0_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_15_io_addInput = mac_1_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_16_clock = clock;
  assign mac_1_16_reset = reset;
  assign mac_1_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_16_io_mulInput = mac_0_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_16_io_addInput = mac_1_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_17_clock = clock;
  assign mac_1_17_reset = reset;
  assign mac_1_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_17_io_mulInput = mac_0_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_17_io_addInput = mac_1_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_18_clock = clock;
  assign mac_1_18_reset = reset;
  assign mac_1_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_18_io_mulInput = mac_0_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_18_io_addInput = mac_1_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_19_clock = clock;
  assign mac_1_19_reset = reset;
  assign mac_1_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_19_io_mulInput = mac_0_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_19_io_addInput = mac_1_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_20_clock = clock;
  assign mac_1_20_reset = reset;
  assign mac_1_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_20_io_mulInput = mac_0_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_20_io_addInput = mac_1_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_21_clock = clock;
  assign mac_1_21_reset = reset;
  assign mac_1_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_21_io_mulInput = mac_0_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_21_io_addInput = mac_1_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_22_clock = clock;
  assign mac_1_22_reset = reset;
  assign mac_1_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_22_io_mulInput = mac_0_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_22_io_addInput = mac_1_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_23_clock = clock;
  assign mac_1_23_reset = reset;
  assign mac_1_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_23_io_mulInput = mac_0_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_23_io_addInput = mac_1_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_24_clock = clock;
  assign mac_1_24_reset = reset;
  assign mac_1_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_24_io_mulInput = mac_0_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_24_io_addInput = mac_1_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_25_clock = clock;
  assign mac_1_25_reset = reset;
  assign mac_1_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_25_io_mulInput = mac_0_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_25_io_addInput = mac_1_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_26_clock = clock;
  assign mac_1_26_reset = reset;
  assign mac_1_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_26_io_mulInput = mac_0_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_26_io_addInput = mac_1_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_27_clock = clock;
  assign mac_1_27_reset = reset;
  assign mac_1_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_27_io_mulInput = mac_0_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_27_io_addInput = mac_1_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_28_clock = clock;
  assign mac_1_28_reset = reset;
  assign mac_1_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_28_io_mulInput = mac_0_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_28_io_addInput = mac_1_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_29_clock = clock;
  assign mac_1_29_reset = reset;
  assign mac_1_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_29_io_mulInput = mac_0_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_29_io_addInput = mac_1_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_30_clock = clock;
  assign mac_1_30_reset = reset;
  assign mac_1_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_30_io_mulInput = mac_0_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_30_io_addInput = mac_1_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_1_31_clock = clock;
  assign mac_1_31_reset = reset;
  assign mac_1_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_1_31_io_mulInput = mac_0_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_1_31_io_addInput = mac_1_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_0_clock = clock;
  assign mac_2_0_reset = reset;
  assign mac_2_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_2_0_io_mulInput = mac_1_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_2_0_io_addInput = bias_2; // @[InnerSystolicArray.scala 57:27]
  assign mac_2_1_clock = clock;
  assign mac_2_1_reset = reset;
  assign mac_2_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_1_io_mulInput = mac_1_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_1_io_addInput = mac_2_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_2_clock = clock;
  assign mac_2_2_reset = reset;
  assign mac_2_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_2_io_mulInput = mac_1_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_2_io_addInput = mac_2_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_3_clock = clock;
  assign mac_2_3_reset = reset;
  assign mac_2_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_3_io_mulInput = mac_1_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_3_io_addInput = mac_2_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_4_clock = clock;
  assign mac_2_4_reset = reset;
  assign mac_2_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_4_io_mulInput = mac_1_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_4_io_addInput = mac_2_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_5_clock = clock;
  assign mac_2_5_reset = reset;
  assign mac_2_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_5_io_mulInput = mac_1_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_5_io_addInput = mac_2_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_6_clock = clock;
  assign mac_2_6_reset = reset;
  assign mac_2_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_6_io_mulInput = mac_1_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_6_io_addInput = mac_2_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_7_clock = clock;
  assign mac_2_7_reset = reset;
  assign mac_2_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_7_io_mulInput = mac_1_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_7_io_addInput = mac_2_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_8_clock = clock;
  assign mac_2_8_reset = reset;
  assign mac_2_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_8_io_mulInput = mac_1_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_8_io_addInput = mac_2_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_9_clock = clock;
  assign mac_2_9_reset = reset;
  assign mac_2_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_9_io_mulInput = mac_1_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_9_io_addInput = mac_2_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_10_clock = clock;
  assign mac_2_10_reset = reset;
  assign mac_2_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_10_io_mulInput = mac_1_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_10_io_addInput = mac_2_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_11_clock = clock;
  assign mac_2_11_reset = reset;
  assign mac_2_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_11_io_mulInput = mac_1_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_11_io_addInput = mac_2_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_12_clock = clock;
  assign mac_2_12_reset = reset;
  assign mac_2_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_12_io_mulInput = mac_1_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_12_io_addInput = mac_2_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_13_clock = clock;
  assign mac_2_13_reset = reset;
  assign mac_2_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_13_io_mulInput = mac_1_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_13_io_addInput = mac_2_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_14_clock = clock;
  assign mac_2_14_reset = reset;
  assign mac_2_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_14_io_mulInput = mac_1_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_14_io_addInput = mac_2_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_15_clock = clock;
  assign mac_2_15_reset = reset;
  assign mac_2_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_15_io_mulInput = mac_1_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_15_io_addInput = mac_2_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_16_clock = clock;
  assign mac_2_16_reset = reset;
  assign mac_2_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_16_io_mulInput = mac_1_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_16_io_addInput = mac_2_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_17_clock = clock;
  assign mac_2_17_reset = reset;
  assign mac_2_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_17_io_mulInput = mac_1_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_17_io_addInput = mac_2_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_18_clock = clock;
  assign mac_2_18_reset = reset;
  assign mac_2_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_18_io_mulInput = mac_1_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_18_io_addInput = mac_2_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_19_clock = clock;
  assign mac_2_19_reset = reset;
  assign mac_2_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_19_io_mulInput = mac_1_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_19_io_addInput = mac_2_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_20_clock = clock;
  assign mac_2_20_reset = reset;
  assign mac_2_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_20_io_mulInput = mac_1_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_20_io_addInput = mac_2_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_21_clock = clock;
  assign mac_2_21_reset = reset;
  assign mac_2_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_21_io_mulInput = mac_1_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_21_io_addInput = mac_2_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_22_clock = clock;
  assign mac_2_22_reset = reset;
  assign mac_2_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_22_io_mulInput = mac_1_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_22_io_addInput = mac_2_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_23_clock = clock;
  assign mac_2_23_reset = reset;
  assign mac_2_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_23_io_mulInput = mac_1_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_23_io_addInput = mac_2_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_24_clock = clock;
  assign mac_2_24_reset = reset;
  assign mac_2_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_24_io_mulInput = mac_1_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_24_io_addInput = mac_2_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_25_clock = clock;
  assign mac_2_25_reset = reset;
  assign mac_2_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_25_io_mulInput = mac_1_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_25_io_addInput = mac_2_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_26_clock = clock;
  assign mac_2_26_reset = reset;
  assign mac_2_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_26_io_mulInput = mac_1_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_26_io_addInput = mac_2_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_27_clock = clock;
  assign mac_2_27_reset = reset;
  assign mac_2_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_27_io_mulInput = mac_1_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_27_io_addInput = mac_2_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_28_clock = clock;
  assign mac_2_28_reset = reset;
  assign mac_2_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_28_io_mulInput = mac_1_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_28_io_addInput = mac_2_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_29_clock = clock;
  assign mac_2_29_reset = reset;
  assign mac_2_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_29_io_mulInput = mac_1_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_29_io_addInput = mac_2_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_30_clock = clock;
  assign mac_2_30_reset = reset;
  assign mac_2_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_30_io_mulInput = mac_1_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_30_io_addInput = mac_2_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_2_31_clock = clock;
  assign mac_2_31_reset = reset;
  assign mac_2_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_2_31_io_mulInput = mac_1_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_2_31_io_addInput = mac_2_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_0_clock = clock;
  assign mac_3_0_reset = reset;
  assign mac_3_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_3_0_io_mulInput = mac_2_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_3_0_io_addInput = bias_3; // @[InnerSystolicArray.scala 57:27]
  assign mac_3_1_clock = clock;
  assign mac_3_1_reset = reset;
  assign mac_3_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_1_io_mulInput = mac_2_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_1_io_addInput = mac_3_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_2_clock = clock;
  assign mac_3_2_reset = reset;
  assign mac_3_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_2_io_mulInput = mac_2_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_2_io_addInput = mac_3_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_3_clock = clock;
  assign mac_3_3_reset = reset;
  assign mac_3_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_3_io_mulInput = mac_2_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_3_io_addInput = mac_3_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_4_clock = clock;
  assign mac_3_4_reset = reset;
  assign mac_3_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_4_io_mulInput = mac_2_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_4_io_addInput = mac_3_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_5_clock = clock;
  assign mac_3_5_reset = reset;
  assign mac_3_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_5_io_mulInput = mac_2_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_5_io_addInput = mac_3_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_6_clock = clock;
  assign mac_3_6_reset = reset;
  assign mac_3_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_6_io_mulInput = mac_2_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_6_io_addInput = mac_3_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_7_clock = clock;
  assign mac_3_7_reset = reset;
  assign mac_3_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_7_io_mulInput = mac_2_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_7_io_addInput = mac_3_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_8_clock = clock;
  assign mac_3_8_reset = reset;
  assign mac_3_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_8_io_mulInput = mac_2_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_8_io_addInput = mac_3_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_9_clock = clock;
  assign mac_3_9_reset = reset;
  assign mac_3_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_9_io_mulInput = mac_2_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_9_io_addInput = mac_3_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_10_clock = clock;
  assign mac_3_10_reset = reset;
  assign mac_3_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_10_io_mulInput = mac_2_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_10_io_addInput = mac_3_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_11_clock = clock;
  assign mac_3_11_reset = reset;
  assign mac_3_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_11_io_mulInput = mac_2_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_11_io_addInput = mac_3_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_12_clock = clock;
  assign mac_3_12_reset = reset;
  assign mac_3_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_12_io_mulInput = mac_2_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_12_io_addInput = mac_3_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_13_clock = clock;
  assign mac_3_13_reset = reset;
  assign mac_3_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_13_io_mulInput = mac_2_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_13_io_addInput = mac_3_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_14_clock = clock;
  assign mac_3_14_reset = reset;
  assign mac_3_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_14_io_mulInput = mac_2_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_14_io_addInput = mac_3_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_15_clock = clock;
  assign mac_3_15_reset = reset;
  assign mac_3_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_15_io_mulInput = mac_2_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_15_io_addInput = mac_3_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_16_clock = clock;
  assign mac_3_16_reset = reset;
  assign mac_3_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_16_io_mulInput = mac_2_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_16_io_addInput = mac_3_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_17_clock = clock;
  assign mac_3_17_reset = reset;
  assign mac_3_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_17_io_mulInput = mac_2_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_17_io_addInput = mac_3_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_18_clock = clock;
  assign mac_3_18_reset = reset;
  assign mac_3_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_18_io_mulInput = mac_2_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_18_io_addInput = mac_3_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_19_clock = clock;
  assign mac_3_19_reset = reset;
  assign mac_3_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_19_io_mulInput = mac_2_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_19_io_addInput = mac_3_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_20_clock = clock;
  assign mac_3_20_reset = reset;
  assign mac_3_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_20_io_mulInput = mac_2_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_20_io_addInput = mac_3_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_21_clock = clock;
  assign mac_3_21_reset = reset;
  assign mac_3_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_21_io_mulInput = mac_2_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_21_io_addInput = mac_3_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_22_clock = clock;
  assign mac_3_22_reset = reset;
  assign mac_3_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_22_io_mulInput = mac_2_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_22_io_addInput = mac_3_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_23_clock = clock;
  assign mac_3_23_reset = reset;
  assign mac_3_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_23_io_mulInput = mac_2_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_23_io_addInput = mac_3_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_24_clock = clock;
  assign mac_3_24_reset = reset;
  assign mac_3_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_24_io_mulInput = mac_2_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_24_io_addInput = mac_3_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_25_clock = clock;
  assign mac_3_25_reset = reset;
  assign mac_3_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_25_io_mulInput = mac_2_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_25_io_addInput = mac_3_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_26_clock = clock;
  assign mac_3_26_reset = reset;
  assign mac_3_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_26_io_mulInput = mac_2_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_26_io_addInput = mac_3_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_27_clock = clock;
  assign mac_3_27_reset = reset;
  assign mac_3_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_27_io_mulInput = mac_2_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_27_io_addInput = mac_3_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_28_clock = clock;
  assign mac_3_28_reset = reset;
  assign mac_3_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_28_io_mulInput = mac_2_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_28_io_addInput = mac_3_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_29_clock = clock;
  assign mac_3_29_reset = reset;
  assign mac_3_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_29_io_mulInput = mac_2_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_29_io_addInput = mac_3_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_30_clock = clock;
  assign mac_3_30_reset = reset;
  assign mac_3_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_30_io_mulInput = mac_2_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_30_io_addInput = mac_3_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_3_31_clock = clock;
  assign mac_3_31_reset = reset;
  assign mac_3_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_3_31_io_mulInput = mac_2_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_3_31_io_addInput = mac_3_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_0_clock = clock;
  assign mac_4_0_reset = reset;
  assign mac_4_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_4_0_io_mulInput = mac_3_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_4_0_io_addInput = bias_4; // @[InnerSystolicArray.scala 57:27]
  assign mac_4_1_clock = clock;
  assign mac_4_1_reset = reset;
  assign mac_4_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_1_io_mulInput = mac_3_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_1_io_addInput = mac_4_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_2_clock = clock;
  assign mac_4_2_reset = reset;
  assign mac_4_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_2_io_mulInput = mac_3_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_2_io_addInput = mac_4_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_3_clock = clock;
  assign mac_4_3_reset = reset;
  assign mac_4_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_3_io_mulInput = mac_3_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_3_io_addInput = mac_4_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_4_clock = clock;
  assign mac_4_4_reset = reset;
  assign mac_4_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_4_io_mulInput = mac_3_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_4_io_addInput = mac_4_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_5_clock = clock;
  assign mac_4_5_reset = reset;
  assign mac_4_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_5_io_mulInput = mac_3_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_5_io_addInput = mac_4_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_6_clock = clock;
  assign mac_4_6_reset = reset;
  assign mac_4_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_6_io_mulInput = mac_3_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_6_io_addInput = mac_4_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_7_clock = clock;
  assign mac_4_7_reset = reset;
  assign mac_4_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_7_io_mulInput = mac_3_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_7_io_addInput = mac_4_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_8_clock = clock;
  assign mac_4_8_reset = reset;
  assign mac_4_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_8_io_mulInput = mac_3_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_8_io_addInput = mac_4_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_9_clock = clock;
  assign mac_4_9_reset = reset;
  assign mac_4_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_9_io_mulInput = mac_3_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_9_io_addInput = mac_4_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_10_clock = clock;
  assign mac_4_10_reset = reset;
  assign mac_4_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_10_io_mulInput = mac_3_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_10_io_addInput = mac_4_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_11_clock = clock;
  assign mac_4_11_reset = reset;
  assign mac_4_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_11_io_mulInput = mac_3_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_11_io_addInput = mac_4_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_12_clock = clock;
  assign mac_4_12_reset = reset;
  assign mac_4_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_12_io_mulInput = mac_3_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_12_io_addInput = mac_4_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_13_clock = clock;
  assign mac_4_13_reset = reset;
  assign mac_4_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_13_io_mulInput = mac_3_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_13_io_addInput = mac_4_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_14_clock = clock;
  assign mac_4_14_reset = reset;
  assign mac_4_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_14_io_mulInput = mac_3_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_14_io_addInput = mac_4_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_15_clock = clock;
  assign mac_4_15_reset = reset;
  assign mac_4_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_15_io_mulInput = mac_3_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_15_io_addInput = mac_4_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_16_clock = clock;
  assign mac_4_16_reset = reset;
  assign mac_4_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_16_io_mulInput = mac_3_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_16_io_addInput = mac_4_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_17_clock = clock;
  assign mac_4_17_reset = reset;
  assign mac_4_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_17_io_mulInput = mac_3_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_17_io_addInput = mac_4_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_18_clock = clock;
  assign mac_4_18_reset = reset;
  assign mac_4_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_18_io_mulInput = mac_3_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_18_io_addInput = mac_4_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_19_clock = clock;
  assign mac_4_19_reset = reset;
  assign mac_4_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_19_io_mulInput = mac_3_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_19_io_addInput = mac_4_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_20_clock = clock;
  assign mac_4_20_reset = reset;
  assign mac_4_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_20_io_mulInput = mac_3_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_20_io_addInput = mac_4_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_21_clock = clock;
  assign mac_4_21_reset = reset;
  assign mac_4_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_21_io_mulInput = mac_3_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_21_io_addInput = mac_4_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_22_clock = clock;
  assign mac_4_22_reset = reset;
  assign mac_4_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_22_io_mulInput = mac_3_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_22_io_addInput = mac_4_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_23_clock = clock;
  assign mac_4_23_reset = reset;
  assign mac_4_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_23_io_mulInput = mac_3_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_23_io_addInput = mac_4_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_24_clock = clock;
  assign mac_4_24_reset = reset;
  assign mac_4_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_24_io_mulInput = mac_3_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_24_io_addInput = mac_4_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_25_clock = clock;
  assign mac_4_25_reset = reset;
  assign mac_4_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_25_io_mulInput = mac_3_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_25_io_addInput = mac_4_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_26_clock = clock;
  assign mac_4_26_reset = reset;
  assign mac_4_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_26_io_mulInput = mac_3_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_26_io_addInput = mac_4_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_27_clock = clock;
  assign mac_4_27_reset = reset;
  assign mac_4_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_27_io_mulInput = mac_3_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_27_io_addInput = mac_4_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_28_clock = clock;
  assign mac_4_28_reset = reset;
  assign mac_4_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_28_io_mulInput = mac_3_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_28_io_addInput = mac_4_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_29_clock = clock;
  assign mac_4_29_reset = reset;
  assign mac_4_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_29_io_mulInput = mac_3_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_29_io_addInput = mac_4_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_30_clock = clock;
  assign mac_4_30_reset = reset;
  assign mac_4_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_30_io_mulInput = mac_3_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_30_io_addInput = mac_4_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_4_31_clock = clock;
  assign mac_4_31_reset = reset;
  assign mac_4_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_4_31_io_mulInput = mac_3_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_4_31_io_addInput = mac_4_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_0_clock = clock;
  assign mac_5_0_reset = reset;
  assign mac_5_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_5_0_io_mulInput = mac_4_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_5_0_io_addInput = bias_5; // @[InnerSystolicArray.scala 57:27]
  assign mac_5_1_clock = clock;
  assign mac_5_1_reset = reset;
  assign mac_5_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_1_io_mulInput = mac_4_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_1_io_addInput = mac_5_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_2_clock = clock;
  assign mac_5_2_reset = reset;
  assign mac_5_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_2_io_mulInput = mac_4_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_2_io_addInput = mac_5_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_3_clock = clock;
  assign mac_5_3_reset = reset;
  assign mac_5_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_3_io_mulInput = mac_4_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_3_io_addInput = mac_5_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_4_clock = clock;
  assign mac_5_4_reset = reset;
  assign mac_5_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_4_io_mulInput = mac_4_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_4_io_addInput = mac_5_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_5_clock = clock;
  assign mac_5_5_reset = reset;
  assign mac_5_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_5_io_mulInput = mac_4_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_5_io_addInput = mac_5_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_6_clock = clock;
  assign mac_5_6_reset = reset;
  assign mac_5_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_6_io_mulInput = mac_4_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_6_io_addInput = mac_5_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_7_clock = clock;
  assign mac_5_7_reset = reset;
  assign mac_5_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_7_io_mulInput = mac_4_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_7_io_addInput = mac_5_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_8_clock = clock;
  assign mac_5_8_reset = reset;
  assign mac_5_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_8_io_mulInput = mac_4_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_8_io_addInput = mac_5_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_9_clock = clock;
  assign mac_5_9_reset = reset;
  assign mac_5_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_9_io_mulInput = mac_4_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_9_io_addInput = mac_5_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_10_clock = clock;
  assign mac_5_10_reset = reset;
  assign mac_5_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_10_io_mulInput = mac_4_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_10_io_addInput = mac_5_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_11_clock = clock;
  assign mac_5_11_reset = reset;
  assign mac_5_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_11_io_mulInput = mac_4_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_11_io_addInput = mac_5_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_12_clock = clock;
  assign mac_5_12_reset = reset;
  assign mac_5_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_12_io_mulInput = mac_4_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_12_io_addInput = mac_5_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_13_clock = clock;
  assign mac_5_13_reset = reset;
  assign mac_5_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_13_io_mulInput = mac_4_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_13_io_addInput = mac_5_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_14_clock = clock;
  assign mac_5_14_reset = reset;
  assign mac_5_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_14_io_mulInput = mac_4_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_14_io_addInput = mac_5_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_15_clock = clock;
  assign mac_5_15_reset = reset;
  assign mac_5_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_15_io_mulInput = mac_4_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_15_io_addInput = mac_5_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_16_clock = clock;
  assign mac_5_16_reset = reset;
  assign mac_5_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_16_io_mulInput = mac_4_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_16_io_addInput = mac_5_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_17_clock = clock;
  assign mac_5_17_reset = reset;
  assign mac_5_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_17_io_mulInput = mac_4_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_17_io_addInput = mac_5_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_18_clock = clock;
  assign mac_5_18_reset = reset;
  assign mac_5_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_18_io_mulInput = mac_4_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_18_io_addInput = mac_5_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_19_clock = clock;
  assign mac_5_19_reset = reset;
  assign mac_5_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_19_io_mulInput = mac_4_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_19_io_addInput = mac_5_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_20_clock = clock;
  assign mac_5_20_reset = reset;
  assign mac_5_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_20_io_mulInput = mac_4_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_20_io_addInput = mac_5_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_21_clock = clock;
  assign mac_5_21_reset = reset;
  assign mac_5_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_21_io_mulInput = mac_4_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_21_io_addInput = mac_5_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_22_clock = clock;
  assign mac_5_22_reset = reset;
  assign mac_5_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_22_io_mulInput = mac_4_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_22_io_addInput = mac_5_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_23_clock = clock;
  assign mac_5_23_reset = reset;
  assign mac_5_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_23_io_mulInput = mac_4_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_23_io_addInput = mac_5_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_24_clock = clock;
  assign mac_5_24_reset = reset;
  assign mac_5_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_24_io_mulInput = mac_4_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_24_io_addInput = mac_5_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_25_clock = clock;
  assign mac_5_25_reset = reset;
  assign mac_5_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_25_io_mulInput = mac_4_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_25_io_addInput = mac_5_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_26_clock = clock;
  assign mac_5_26_reset = reset;
  assign mac_5_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_26_io_mulInput = mac_4_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_26_io_addInput = mac_5_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_27_clock = clock;
  assign mac_5_27_reset = reset;
  assign mac_5_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_27_io_mulInput = mac_4_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_27_io_addInput = mac_5_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_28_clock = clock;
  assign mac_5_28_reset = reset;
  assign mac_5_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_28_io_mulInput = mac_4_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_28_io_addInput = mac_5_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_29_clock = clock;
  assign mac_5_29_reset = reset;
  assign mac_5_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_29_io_mulInput = mac_4_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_29_io_addInput = mac_5_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_30_clock = clock;
  assign mac_5_30_reset = reset;
  assign mac_5_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_30_io_mulInput = mac_4_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_30_io_addInput = mac_5_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_5_31_clock = clock;
  assign mac_5_31_reset = reset;
  assign mac_5_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_5_31_io_mulInput = mac_4_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_5_31_io_addInput = mac_5_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_0_clock = clock;
  assign mac_6_0_reset = reset;
  assign mac_6_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_6_0_io_mulInput = mac_5_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_6_0_io_addInput = bias_6; // @[InnerSystolicArray.scala 57:27]
  assign mac_6_1_clock = clock;
  assign mac_6_1_reset = reset;
  assign mac_6_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_1_io_mulInput = mac_5_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_1_io_addInput = mac_6_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_2_clock = clock;
  assign mac_6_2_reset = reset;
  assign mac_6_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_2_io_mulInput = mac_5_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_2_io_addInput = mac_6_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_3_clock = clock;
  assign mac_6_3_reset = reset;
  assign mac_6_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_3_io_mulInput = mac_5_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_3_io_addInput = mac_6_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_4_clock = clock;
  assign mac_6_4_reset = reset;
  assign mac_6_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_4_io_mulInput = mac_5_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_4_io_addInput = mac_6_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_5_clock = clock;
  assign mac_6_5_reset = reset;
  assign mac_6_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_5_io_mulInput = mac_5_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_5_io_addInput = mac_6_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_6_clock = clock;
  assign mac_6_6_reset = reset;
  assign mac_6_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_6_io_mulInput = mac_5_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_6_io_addInput = mac_6_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_7_clock = clock;
  assign mac_6_7_reset = reset;
  assign mac_6_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_7_io_mulInput = mac_5_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_7_io_addInput = mac_6_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_8_clock = clock;
  assign mac_6_8_reset = reset;
  assign mac_6_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_8_io_mulInput = mac_5_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_8_io_addInput = mac_6_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_9_clock = clock;
  assign mac_6_9_reset = reset;
  assign mac_6_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_9_io_mulInput = mac_5_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_9_io_addInput = mac_6_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_10_clock = clock;
  assign mac_6_10_reset = reset;
  assign mac_6_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_10_io_mulInput = mac_5_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_10_io_addInput = mac_6_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_11_clock = clock;
  assign mac_6_11_reset = reset;
  assign mac_6_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_11_io_mulInput = mac_5_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_11_io_addInput = mac_6_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_12_clock = clock;
  assign mac_6_12_reset = reset;
  assign mac_6_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_12_io_mulInput = mac_5_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_12_io_addInput = mac_6_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_13_clock = clock;
  assign mac_6_13_reset = reset;
  assign mac_6_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_13_io_mulInput = mac_5_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_13_io_addInput = mac_6_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_14_clock = clock;
  assign mac_6_14_reset = reset;
  assign mac_6_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_14_io_mulInput = mac_5_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_14_io_addInput = mac_6_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_15_clock = clock;
  assign mac_6_15_reset = reset;
  assign mac_6_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_15_io_mulInput = mac_5_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_15_io_addInput = mac_6_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_16_clock = clock;
  assign mac_6_16_reset = reset;
  assign mac_6_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_16_io_mulInput = mac_5_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_16_io_addInput = mac_6_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_17_clock = clock;
  assign mac_6_17_reset = reset;
  assign mac_6_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_17_io_mulInput = mac_5_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_17_io_addInput = mac_6_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_18_clock = clock;
  assign mac_6_18_reset = reset;
  assign mac_6_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_18_io_mulInput = mac_5_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_18_io_addInput = mac_6_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_19_clock = clock;
  assign mac_6_19_reset = reset;
  assign mac_6_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_19_io_mulInput = mac_5_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_19_io_addInput = mac_6_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_20_clock = clock;
  assign mac_6_20_reset = reset;
  assign mac_6_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_20_io_mulInput = mac_5_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_20_io_addInput = mac_6_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_21_clock = clock;
  assign mac_6_21_reset = reset;
  assign mac_6_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_21_io_mulInput = mac_5_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_21_io_addInput = mac_6_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_22_clock = clock;
  assign mac_6_22_reset = reset;
  assign mac_6_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_22_io_mulInput = mac_5_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_22_io_addInput = mac_6_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_23_clock = clock;
  assign mac_6_23_reset = reset;
  assign mac_6_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_23_io_mulInput = mac_5_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_23_io_addInput = mac_6_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_24_clock = clock;
  assign mac_6_24_reset = reset;
  assign mac_6_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_24_io_mulInput = mac_5_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_24_io_addInput = mac_6_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_25_clock = clock;
  assign mac_6_25_reset = reset;
  assign mac_6_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_25_io_mulInput = mac_5_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_25_io_addInput = mac_6_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_26_clock = clock;
  assign mac_6_26_reset = reset;
  assign mac_6_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_26_io_mulInput = mac_5_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_26_io_addInput = mac_6_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_27_clock = clock;
  assign mac_6_27_reset = reset;
  assign mac_6_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_27_io_mulInput = mac_5_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_27_io_addInput = mac_6_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_28_clock = clock;
  assign mac_6_28_reset = reset;
  assign mac_6_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_28_io_mulInput = mac_5_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_28_io_addInput = mac_6_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_29_clock = clock;
  assign mac_6_29_reset = reset;
  assign mac_6_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_29_io_mulInput = mac_5_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_29_io_addInput = mac_6_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_30_clock = clock;
  assign mac_6_30_reset = reset;
  assign mac_6_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_30_io_mulInput = mac_5_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_30_io_addInput = mac_6_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_6_31_clock = clock;
  assign mac_6_31_reset = reset;
  assign mac_6_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_6_31_io_mulInput = mac_5_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_6_31_io_addInput = mac_6_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_0_clock = clock;
  assign mac_7_0_reset = reset;
  assign mac_7_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_7_0_io_mulInput = mac_6_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_7_0_io_addInput = bias_7; // @[InnerSystolicArray.scala 57:27]
  assign mac_7_1_clock = clock;
  assign mac_7_1_reset = reset;
  assign mac_7_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_1_io_mulInput = mac_6_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_1_io_addInput = mac_7_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_2_clock = clock;
  assign mac_7_2_reset = reset;
  assign mac_7_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_2_io_mulInput = mac_6_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_2_io_addInput = mac_7_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_3_clock = clock;
  assign mac_7_3_reset = reset;
  assign mac_7_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_3_io_mulInput = mac_6_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_3_io_addInput = mac_7_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_4_clock = clock;
  assign mac_7_4_reset = reset;
  assign mac_7_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_4_io_mulInput = mac_6_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_4_io_addInput = mac_7_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_5_clock = clock;
  assign mac_7_5_reset = reset;
  assign mac_7_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_5_io_mulInput = mac_6_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_5_io_addInput = mac_7_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_6_clock = clock;
  assign mac_7_6_reset = reset;
  assign mac_7_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_6_io_mulInput = mac_6_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_6_io_addInput = mac_7_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_7_clock = clock;
  assign mac_7_7_reset = reset;
  assign mac_7_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_7_io_mulInput = mac_6_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_7_io_addInput = mac_7_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_8_clock = clock;
  assign mac_7_8_reset = reset;
  assign mac_7_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_8_io_mulInput = mac_6_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_8_io_addInput = mac_7_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_9_clock = clock;
  assign mac_7_9_reset = reset;
  assign mac_7_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_9_io_mulInput = mac_6_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_9_io_addInput = mac_7_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_10_clock = clock;
  assign mac_7_10_reset = reset;
  assign mac_7_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_10_io_mulInput = mac_6_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_10_io_addInput = mac_7_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_11_clock = clock;
  assign mac_7_11_reset = reset;
  assign mac_7_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_11_io_mulInput = mac_6_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_11_io_addInput = mac_7_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_12_clock = clock;
  assign mac_7_12_reset = reset;
  assign mac_7_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_12_io_mulInput = mac_6_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_12_io_addInput = mac_7_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_13_clock = clock;
  assign mac_7_13_reset = reset;
  assign mac_7_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_13_io_mulInput = mac_6_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_13_io_addInput = mac_7_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_14_clock = clock;
  assign mac_7_14_reset = reset;
  assign mac_7_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_14_io_mulInput = mac_6_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_14_io_addInput = mac_7_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_15_clock = clock;
  assign mac_7_15_reset = reset;
  assign mac_7_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_15_io_mulInput = mac_6_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_15_io_addInput = mac_7_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_16_clock = clock;
  assign mac_7_16_reset = reset;
  assign mac_7_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_16_io_mulInput = mac_6_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_16_io_addInput = mac_7_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_17_clock = clock;
  assign mac_7_17_reset = reset;
  assign mac_7_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_17_io_mulInput = mac_6_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_17_io_addInput = mac_7_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_18_clock = clock;
  assign mac_7_18_reset = reset;
  assign mac_7_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_18_io_mulInput = mac_6_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_18_io_addInput = mac_7_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_19_clock = clock;
  assign mac_7_19_reset = reset;
  assign mac_7_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_19_io_mulInput = mac_6_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_19_io_addInput = mac_7_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_20_clock = clock;
  assign mac_7_20_reset = reset;
  assign mac_7_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_20_io_mulInput = mac_6_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_20_io_addInput = mac_7_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_21_clock = clock;
  assign mac_7_21_reset = reset;
  assign mac_7_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_21_io_mulInput = mac_6_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_21_io_addInput = mac_7_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_22_clock = clock;
  assign mac_7_22_reset = reset;
  assign mac_7_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_22_io_mulInput = mac_6_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_22_io_addInput = mac_7_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_23_clock = clock;
  assign mac_7_23_reset = reset;
  assign mac_7_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_23_io_mulInput = mac_6_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_23_io_addInput = mac_7_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_24_clock = clock;
  assign mac_7_24_reset = reset;
  assign mac_7_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_24_io_mulInput = mac_6_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_24_io_addInput = mac_7_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_25_clock = clock;
  assign mac_7_25_reset = reset;
  assign mac_7_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_25_io_mulInput = mac_6_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_25_io_addInput = mac_7_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_26_clock = clock;
  assign mac_7_26_reset = reset;
  assign mac_7_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_26_io_mulInput = mac_6_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_26_io_addInput = mac_7_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_27_clock = clock;
  assign mac_7_27_reset = reset;
  assign mac_7_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_27_io_mulInput = mac_6_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_27_io_addInput = mac_7_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_28_clock = clock;
  assign mac_7_28_reset = reset;
  assign mac_7_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_28_io_mulInput = mac_6_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_28_io_addInput = mac_7_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_29_clock = clock;
  assign mac_7_29_reset = reset;
  assign mac_7_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_29_io_mulInput = mac_6_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_29_io_addInput = mac_7_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_30_clock = clock;
  assign mac_7_30_reset = reset;
  assign mac_7_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_30_io_mulInput = mac_6_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_30_io_addInput = mac_7_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_7_31_clock = clock;
  assign mac_7_31_reset = reset;
  assign mac_7_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_7_31_io_mulInput = mac_6_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_7_31_io_addInput = mac_7_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_0_clock = clock;
  assign mac_8_0_reset = reset;
  assign mac_8_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_8_0_io_mulInput = mac_7_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_8_0_io_addInput = bias_8; // @[InnerSystolicArray.scala 57:27]
  assign mac_8_1_clock = clock;
  assign mac_8_1_reset = reset;
  assign mac_8_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_1_io_mulInput = mac_7_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_1_io_addInput = mac_8_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_2_clock = clock;
  assign mac_8_2_reset = reset;
  assign mac_8_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_2_io_mulInput = mac_7_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_2_io_addInput = mac_8_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_3_clock = clock;
  assign mac_8_3_reset = reset;
  assign mac_8_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_3_io_mulInput = mac_7_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_3_io_addInput = mac_8_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_4_clock = clock;
  assign mac_8_4_reset = reset;
  assign mac_8_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_4_io_mulInput = mac_7_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_4_io_addInput = mac_8_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_5_clock = clock;
  assign mac_8_5_reset = reset;
  assign mac_8_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_5_io_mulInput = mac_7_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_5_io_addInput = mac_8_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_6_clock = clock;
  assign mac_8_6_reset = reset;
  assign mac_8_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_6_io_mulInput = mac_7_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_6_io_addInput = mac_8_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_7_clock = clock;
  assign mac_8_7_reset = reset;
  assign mac_8_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_7_io_mulInput = mac_7_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_7_io_addInput = mac_8_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_8_clock = clock;
  assign mac_8_8_reset = reset;
  assign mac_8_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_8_io_mulInput = mac_7_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_8_io_addInput = mac_8_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_9_clock = clock;
  assign mac_8_9_reset = reset;
  assign mac_8_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_9_io_mulInput = mac_7_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_9_io_addInput = mac_8_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_10_clock = clock;
  assign mac_8_10_reset = reset;
  assign mac_8_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_10_io_mulInput = mac_7_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_10_io_addInput = mac_8_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_11_clock = clock;
  assign mac_8_11_reset = reset;
  assign mac_8_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_11_io_mulInput = mac_7_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_11_io_addInput = mac_8_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_12_clock = clock;
  assign mac_8_12_reset = reset;
  assign mac_8_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_12_io_mulInput = mac_7_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_12_io_addInput = mac_8_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_13_clock = clock;
  assign mac_8_13_reset = reset;
  assign mac_8_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_13_io_mulInput = mac_7_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_13_io_addInput = mac_8_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_14_clock = clock;
  assign mac_8_14_reset = reset;
  assign mac_8_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_14_io_mulInput = mac_7_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_14_io_addInput = mac_8_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_15_clock = clock;
  assign mac_8_15_reset = reset;
  assign mac_8_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_15_io_mulInput = mac_7_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_15_io_addInput = mac_8_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_16_clock = clock;
  assign mac_8_16_reset = reset;
  assign mac_8_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_16_io_mulInput = mac_7_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_16_io_addInput = mac_8_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_17_clock = clock;
  assign mac_8_17_reset = reset;
  assign mac_8_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_17_io_mulInput = mac_7_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_17_io_addInput = mac_8_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_18_clock = clock;
  assign mac_8_18_reset = reset;
  assign mac_8_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_18_io_mulInput = mac_7_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_18_io_addInput = mac_8_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_19_clock = clock;
  assign mac_8_19_reset = reset;
  assign mac_8_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_19_io_mulInput = mac_7_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_19_io_addInput = mac_8_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_20_clock = clock;
  assign mac_8_20_reset = reset;
  assign mac_8_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_20_io_mulInput = mac_7_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_20_io_addInput = mac_8_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_21_clock = clock;
  assign mac_8_21_reset = reset;
  assign mac_8_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_21_io_mulInput = mac_7_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_21_io_addInput = mac_8_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_22_clock = clock;
  assign mac_8_22_reset = reset;
  assign mac_8_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_22_io_mulInput = mac_7_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_22_io_addInput = mac_8_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_23_clock = clock;
  assign mac_8_23_reset = reset;
  assign mac_8_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_23_io_mulInput = mac_7_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_23_io_addInput = mac_8_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_24_clock = clock;
  assign mac_8_24_reset = reset;
  assign mac_8_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_24_io_mulInput = mac_7_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_24_io_addInput = mac_8_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_25_clock = clock;
  assign mac_8_25_reset = reset;
  assign mac_8_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_25_io_mulInput = mac_7_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_25_io_addInput = mac_8_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_26_clock = clock;
  assign mac_8_26_reset = reset;
  assign mac_8_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_26_io_mulInput = mac_7_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_26_io_addInput = mac_8_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_27_clock = clock;
  assign mac_8_27_reset = reset;
  assign mac_8_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_27_io_mulInput = mac_7_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_27_io_addInput = mac_8_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_28_clock = clock;
  assign mac_8_28_reset = reset;
  assign mac_8_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_28_io_mulInput = mac_7_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_28_io_addInput = mac_8_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_29_clock = clock;
  assign mac_8_29_reset = reset;
  assign mac_8_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_29_io_mulInput = mac_7_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_29_io_addInput = mac_8_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_30_clock = clock;
  assign mac_8_30_reset = reset;
  assign mac_8_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_30_io_mulInput = mac_7_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_30_io_addInput = mac_8_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_8_31_clock = clock;
  assign mac_8_31_reset = reset;
  assign mac_8_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_8_31_io_mulInput = mac_7_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_8_31_io_addInput = mac_8_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_0_clock = clock;
  assign mac_9_0_reset = reset;
  assign mac_9_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_9_0_io_mulInput = mac_8_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_9_0_io_addInput = bias_9; // @[InnerSystolicArray.scala 57:27]
  assign mac_9_1_clock = clock;
  assign mac_9_1_reset = reset;
  assign mac_9_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_1_io_mulInput = mac_8_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_1_io_addInput = mac_9_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_2_clock = clock;
  assign mac_9_2_reset = reset;
  assign mac_9_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_2_io_mulInput = mac_8_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_2_io_addInput = mac_9_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_3_clock = clock;
  assign mac_9_3_reset = reset;
  assign mac_9_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_3_io_mulInput = mac_8_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_3_io_addInput = mac_9_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_4_clock = clock;
  assign mac_9_4_reset = reset;
  assign mac_9_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_4_io_mulInput = mac_8_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_4_io_addInput = mac_9_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_5_clock = clock;
  assign mac_9_5_reset = reset;
  assign mac_9_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_5_io_mulInput = mac_8_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_5_io_addInput = mac_9_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_6_clock = clock;
  assign mac_9_6_reset = reset;
  assign mac_9_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_6_io_mulInput = mac_8_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_6_io_addInput = mac_9_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_7_clock = clock;
  assign mac_9_7_reset = reset;
  assign mac_9_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_7_io_mulInput = mac_8_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_7_io_addInput = mac_9_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_8_clock = clock;
  assign mac_9_8_reset = reset;
  assign mac_9_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_8_io_mulInput = mac_8_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_8_io_addInput = mac_9_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_9_clock = clock;
  assign mac_9_9_reset = reset;
  assign mac_9_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_9_io_mulInput = mac_8_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_9_io_addInput = mac_9_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_10_clock = clock;
  assign mac_9_10_reset = reset;
  assign mac_9_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_10_io_mulInput = mac_8_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_10_io_addInput = mac_9_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_11_clock = clock;
  assign mac_9_11_reset = reset;
  assign mac_9_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_11_io_mulInput = mac_8_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_11_io_addInput = mac_9_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_12_clock = clock;
  assign mac_9_12_reset = reset;
  assign mac_9_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_12_io_mulInput = mac_8_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_12_io_addInput = mac_9_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_13_clock = clock;
  assign mac_9_13_reset = reset;
  assign mac_9_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_13_io_mulInput = mac_8_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_13_io_addInput = mac_9_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_14_clock = clock;
  assign mac_9_14_reset = reset;
  assign mac_9_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_14_io_mulInput = mac_8_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_14_io_addInput = mac_9_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_15_clock = clock;
  assign mac_9_15_reset = reset;
  assign mac_9_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_15_io_mulInput = mac_8_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_15_io_addInput = mac_9_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_16_clock = clock;
  assign mac_9_16_reset = reset;
  assign mac_9_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_16_io_mulInput = mac_8_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_16_io_addInput = mac_9_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_17_clock = clock;
  assign mac_9_17_reset = reset;
  assign mac_9_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_17_io_mulInput = mac_8_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_17_io_addInput = mac_9_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_18_clock = clock;
  assign mac_9_18_reset = reset;
  assign mac_9_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_18_io_mulInput = mac_8_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_18_io_addInput = mac_9_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_19_clock = clock;
  assign mac_9_19_reset = reset;
  assign mac_9_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_19_io_mulInput = mac_8_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_19_io_addInput = mac_9_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_20_clock = clock;
  assign mac_9_20_reset = reset;
  assign mac_9_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_20_io_mulInput = mac_8_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_20_io_addInput = mac_9_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_21_clock = clock;
  assign mac_9_21_reset = reset;
  assign mac_9_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_21_io_mulInput = mac_8_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_21_io_addInput = mac_9_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_22_clock = clock;
  assign mac_9_22_reset = reset;
  assign mac_9_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_22_io_mulInput = mac_8_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_22_io_addInput = mac_9_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_23_clock = clock;
  assign mac_9_23_reset = reset;
  assign mac_9_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_23_io_mulInput = mac_8_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_23_io_addInput = mac_9_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_24_clock = clock;
  assign mac_9_24_reset = reset;
  assign mac_9_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_24_io_mulInput = mac_8_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_24_io_addInput = mac_9_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_25_clock = clock;
  assign mac_9_25_reset = reset;
  assign mac_9_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_25_io_mulInput = mac_8_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_25_io_addInput = mac_9_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_26_clock = clock;
  assign mac_9_26_reset = reset;
  assign mac_9_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_26_io_mulInput = mac_8_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_26_io_addInput = mac_9_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_27_clock = clock;
  assign mac_9_27_reset = reset;
  assign mac_9_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_27_io_mulInput = mac_8_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_27_io_addInput = mac_9_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_28_clock = clock;
  assign mac_9_28_reset = reset;
  assign mac_9_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_28_io_mulInput = mac_8_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_28_io_addInput = mac_9_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_29_clock = clock;
  assign mac_9_29_reset = reset;
  assign mac_9_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_29_io_mulInput = mac_8_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_29_io_addInput = mac_9_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_30_clock = clock;
  assign mac_9_30_reset = reset;
  assign mac_9_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_30_io_mulInput = mac_8_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_30_io_addInput = mac_9_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_9_31_clock = clock;
  assign mac_9_31_reset = reset;
  assign mac_9_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_9_31_io_mulInput = mac_8_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_9_31_io_addInput = mac_9_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_0_clock = clock;
  assign mac_10_0_reset = reset;
  assign mac_10_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_10_0_io_mulInput = mac_9_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_10_0_io_addInput = bias_10; // @[InnerSystolicArray.scala 57:27]
  assign mac_10_1_clock = clock;
  assign mac_10_1_reset = reset;
  assign mac_10_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_1_io_mulInput = mac_9_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_1_io_addInput = mac_10_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_2_clock = clock;
  assign mac_10_2_reset = reset;
  assign mac_10_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_2_io_mulInput = mac_9_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_2_io_addInput = mac_10_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_3_clock = clock;
  assign mac_10_3_reset = reset;
  assign mac_10_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_3_io_mulInput = mac_9_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_3_io_addInput = mac_10_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_4_clock = clock;
  assign mac_10_4_reset = reset;
  assign mac_10_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_4_io_mulInput = mac_9_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_4_io_addInput = mac_10_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_5_clock = clock;
  assign mac_10_5_reset = reset;
  assign mac_10_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_5_io_mulInput = mac_9_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_5_io_addInput = mac_10_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_6_clock = clock;
  assign mac_10_6_reset = reset;
  assign mac_10_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_6_io_mulInput = mac_9_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_6_io_addInput = mac_10_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_7_clock = clock;
  assign mac_10_7_reset = reset;
  assign mac_10_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_7_io_mulInput = mac_9_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_7_io_addInput = mac_10_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_8_clock = clock;
  assign mac_10_8_reset = reset;
  assign mac_10_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_8_io_mulInput = mac_9_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_8_io_addInput = mac_10_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_9_clock = clock;
  assign mac_10_9_reset = reset;
  assign mac_10_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_9_io_mulInput = mac_9_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_9_io_addInput = mac_10_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_10_clock = clock;
  assign mac_10_10_reset = reset;
  assign mac_10_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_10_io_mulInput = mac_9_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_10_io_addInput = mac_10_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_11_clock = clock;
  assign mac_10_11_reset = reset;
  assign mac_10_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_11_io_mulInput = mac_9_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_11_io_addInput = mac_10_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_12_clock = clock;
  assign mac_10_12_reset = reset;
  assign mac_10_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_12_io_mulInput = mac_9_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_12_io_addInput = mac_10_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_13_clock = clock;
  assign mac_10_13_reset = reset;
  assign mac_10_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_13_io_mulInput = mac_9_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_13_io_addInput = mac_10_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_14_clock = clock;
  assign mac_10_14_reset = reset;
  assign mac_10_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_14_io_mulInput = mac_9_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_14_io_addInput = mac_10_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_15_clock = clock;
  assign mac_10_15_reset = reset;
  assign mac_10_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_15_io_mulInput = mac_9_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_15_io_addInput = mac_10_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_16_clock = clock;
  assign mac_10_16_reset = reset;
  assign mac_10_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_16_io_mulInput = mac_9_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_16_io_addInput = mac_10_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_17_clock = clock;
  assign mac_10_17_reset = reset;
  assign mac_10_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_17_io_mulInput = mac_9_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_17_io_addInput = mac_10_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_18_clock = clock;
  assign mac_10_18_reset = reset;
  assign mac_10_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_18_io_mulInput = mac_9_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_18_io_addInput = mac_10_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_19_clock = clock;
  assign mac_10_19_reset = reset;
  assign mac_10_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_19_io_mulInput = mac_9_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_19_io_addInput = mac_10_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_20_clock = clock;
  assign mac_10_20_reset = reset;
  assign mac_10_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_20_io_mulInput = mac_9_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_20_io_addInput = mac_10_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_21_clock = clock;
  assign mac_10_21_reset = reset;
  assign mac_10_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_21_io_mulInput = mac_9_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_21_io_addInput = mac_10_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_22_clock = clock;
  assign mac_10_22_reset = reset;
  assign mac_10_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_22_io_mulInput = mac_9_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_22_io_addInput = mac_10_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_23_clock = clock;
  assign mac_10_23_reset = reset;
  assign mac_10_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_23_io_mulInput = mac_9_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_23_io_addInput = mac_10_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_24_clock = clock;
  assign mac_10_24_reset = reset;
  assign mac_10_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_24_io_mulInput = mac_9_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_24_io_addInput = mac_10_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_25_clock = clock;
  assign mac_10_25_reset = reset;
  assign mac_10_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_25_io_mulInput = mac_9_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_25_io_addInput = mac_10_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_26_clock = clock;
  assign mac_10_26_reset = reset;
  assign mac_10_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_26_io_mulInput = mac_9_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_26_io_addInput = mac_10_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_27_clock = clock;
  assign mac_10_27_reset = reset;
  assign mac_10_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_27_io_mulInput = mac_9_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_27_io_addInput = mac_10_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_28_clock = clock;
  assign mac_10_28_reset = reset;
  assign mac_10_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_28_io_mulInput = mac_9_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_28_io_addInput = mac_10_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_29_clock = clock;
  assign mac_10_29_reset = reset;
  assign mac_10_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_29_io_mulInput = mac_9_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_29_io_addInput = mac_10_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_30_clock = clock;
  assign mac_10_30_reset = reset;
  assign mac_10_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_30_io_mulInput = mac_9_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_30_io_addInput = mac_10_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_10_31_clock = clock;
  assign mac_10_31_reset = reset;
  assign mac_10_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_10_31_io_mulInput = mac_9_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_10_31_io_addInput = mac_10_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_0_clock = clock;
  assign mac_11_0_reset = reset;
  assign mac_11_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_11_0_io_mulInput = mac_10_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_11_0_io_addInput = bias_11; // @[InnerSystolicArray.scala 57:27]
  assign mac_11_1_clock = clock;
  assign mac_11_1_reset = reset;
  assign mac_11_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_1_io_mulInput = mac_10_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_1_io_addInput = mac_11_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_2_clock = clock;
  assign mac_11_2_reset = reset;
  assign mac_11_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_2_io_mulInput = mac_10_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_2_io_addInput = mac_11_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_3_clock = clock;
  assign mac_11_3_reset = reset;
  assign mac_11_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_3_io_mulInput = mac_10_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_3_io_addInput = mac_11_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_4_clock = clock;
  assign mac_11_4_reset = reset;
  assign mac_11_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_4_io_mulInput = mac_10_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_4_io_addInput = mac_11_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_5_clock = clock;
  assign mac_11_5_reset = reset;
  assign mac_11_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_5_io_mulInput = mac_10_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_5_io_addInput = mac_11_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_6_clock = clock;
  assign mac_11_6_reset = reset;
  assign mac_11_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_6_io_mulInput = mac_10_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_6_io_addInput = mac_11_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_7_clock = clock;
  assign mac_11_7_reset = reset;
  assign mac_11_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_7_io_mulInput = mac_10_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_7_io_addInput = mac_11_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_8_clock = clock;
  assign mac_11_8_reset = reset;
  assign mac_11_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_8_io_mulInput = mac_10_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_8_io_addInput = mac_11_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_9_clock = clock;
  assign mac_11_9_reset = reset;
  assign mac_11_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_9_io_mulInput = mac_10_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_9_io_addInput = mac_11_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_10_clock = clock;
  assign mac_11_10_reset = reset;
  assign mac_11_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_10_io_mulInput = mac_10_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_10_io_addInput = mac_11_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_11_clock = clock;
  assign mac_11_11_reset = reset;
  assign mac_11_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_11_io_mulInput = mac_10_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_11_io_addInput = mac_11_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_12_clock = clock;
  assign mac_11_12_reset = reset;
  assign mac_11_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_12_io_mulInput = mac_10_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_12_io_addInput = mac_11_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_13_clock = clock;
  assign mac_11_13_reset = reset;
  assign mac_11_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_13_io_mulInput = mac_10_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_13_io_addInput = mac_11_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_14_clock = clock;
  assign mac_11_14_reset = reset;
  assign mac_11_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_14_io_mulInput = mac_10_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_14_io_addInput = mac_11_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_15_clock = clock;
  assign mac_11_15_reset = reset;
  assign mac_11_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_15_io_mulInput = mac_10_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_15_io_addInput = mac_11_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_16_clock = clock;
  assign mac_11_16_reset = reset;
  assign mac_11_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_16_io_mulInput = mac_10_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_16_io_addInput = mac_11_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_17_clock = clock;
  assign mac_11_17_reset = reset;
  assign mac_11_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_17_io_mulInput = mac_10_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_17_io_addInput = mac_11_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_18_clock = clock;
  assign mac_11_18_reset = reset;
  assign mac_11_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_18_io_mulInput = mac_10_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_18_io_addInput = mac_11_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_19_clock = clock;
  assign mac_11_19_reset = reset;
  assign mac_11_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_19_io_mulInput = mac_10_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_19_io_addInput = mac_11_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_20_clock = clock;
  assign mac_11_20_reset = reset;
  assign mac_11_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_20_io_mulInput = mac_10_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_20_io_addInput = mac_11_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_21_clock = clock;
  assign mac_11_21_reset = reset;
  assign mac_11_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_21_io_mulInput = mac_10_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_21_io_addInput = mac_11_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_22_clock = clock;
  assign mac_11_22_reset = reset;
  assign mac_11_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_22_io_mulInput = mac_10_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_22_io_addInput = mac_11_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_23_clock = clock;
  assign mac_11_23_reset = reset;
  assign mac_11_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_23_io_mulInput = mac_10_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_23_io_addInput = mac_11_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_24_clock = clock;
  assign mac_11_24_reset = reset;
  assign mac_11_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_24_io_mulInput = mac_10_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_24_io_addInput = mac_11_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_25_clock = clock;
  assign mac_11_25_reset = reset;
  assign mac_11_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_25_io_mulInput = mac_10_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_25_io_addInput = mac_11_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_26_clock = clock;
  assign mac_11_26_reset = reset;
  assign mac_11_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_26_io_mulInput = mac_10_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_26_io_addInput = mac_11_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_27_clock = clock;
  assign mac_11_27_reset = reset;
  assign mac_11_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_27_io_mulInput = mac_10_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_27_io_addInput = mac_11_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_28_clock = clock;
  assign mac_11_28_reset = reset;
  assign mac_11_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_28_io_mulInput = mac_10_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_28_io_addInput = mac_11_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_29_clock = clock;
  assign mac_11_29_reset = reset;
  assign mac_11_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_29_io_mulInput = mac_10_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_29_io_addInput = mac_11_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_30_clock = clock;
  assign mac_11_30_reset = reset;
  assign mac_11_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_30_io_mulInput = mac_10_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_30_io_addInput = mac_11_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_11_31_clock = clock;
  assign mac_11_31_reset = reset;
  assign mac_11_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_11_31_io_mulInput = mac_10_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_11_31_io_addInput = mac_11_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_0_clock = clock;
  assign mac_12_0_reset = reset;
  assign mac_12_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_12_0_io_mulInput = mac_11_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_12_0_io_addInput = bias_12; // @[InnerSystolicArray.scala 57:27]
  assign mac_12_1_clock = clock;
  assign mac_12_1_reset = reset;
  assign mac_12_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_1_io_mulInput = mac_11_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_1_io_addInput = mac_12_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_2_clock = clock;
  assign mac_12_2_reset = reset;
  assign mac_12_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_2_io_mulInput = mac_11_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_2_io_addInput = mac_12_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_3_clock = clock;
  assign mac_12_3_reset = reset;
  assign mac_12_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_3_io_mulInput = mac_11_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_3_io_addInput = mac_12_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_4_clock = clock;
  assign mac_12_4_reset = reset;
  assign mac_12_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_4_io_mulInput = mac_11_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_4_io_addInput = mac_12_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_5_clock = clock;
  assign mac_12_5_reset = reset;
  assign mac_12_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_5_io_mulInput = mac_11_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_5_io_addInput = mac_12_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_6_clock = clock;
  assign mac_12_6_reset = reset;
  assign mac_12_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_6_io_mulInput = mac_11_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_6_io_addInput = mac_12_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_7_clock = clock;
  assign mac_12_7_reset = reset;
  assign mac_12_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_7_io_mulInput = mac_11_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_7_io_addInput = mac_12_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_8_clock = clock;
  assign mac_12_8_reset = reset;
  assign mac_12_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_8_io_mulInput = mac_11_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_8_io_addInput = mac_12_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_9_clock = clock;
  assign mac_12_9_reset = reset;
  assign mac_12_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_9_io_mulInput = mac_11_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_9_io_addInput = mac_12_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_10_clock = clock;
  assign mac_12_10_reset = reset;
  assign mac_12_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_10_io_mulInput = mac_11_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_10_io_addInput = mac_12_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_11_clock = clock;
  assign mac_12_11_reset = reset;
  assign mac_12_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_11_io_mulInput = mac_11_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_11_io_addInput = mac_12_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_12_clock = clock;
  assign mac_12_12_reset = reset;
  assign mac_12_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_12_io_mulInput = mac_11_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_12_io_addInput = mac_12_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_13_clock = clock;
  assign mac_12_13_reset = reset;
  assign mac_12_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_13_io_mulInput = mac_11_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_13_io_addInput = mac_12_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_14_clock = clock;
  assign mac_12_14_reset = reset;
  assign mac_12_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_14_io_mulInput = mac_11_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_14_io_addInput = mac_12_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_15_clock = clock;
  assign mac_12_15_reset = reset;
  assign mac_12_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_15_io_mulInput = mac_11_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_15_io_addInput = mac_12_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_16_clock = clock;
  assign mac_12_16_reset = reset;
  assign mac_12_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_16_io_mulInput = mac_11_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_16_io_addInput = mac_12_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_17_clock = clock;
  assign mac_12_17_reset = reset;
  assign mac_12_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_17_io_mulInput = mac_11_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_17_io_addInput = mac_12_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_18_clock = clock;
  assign mac_12_18_reset = reset;
  assign mac_12_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_18_io_mulInput = mac_11_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_18_io_addInput = mac_12_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_19_clock = clock;
  assign mac_12_19_reset = reset;
  assign mac_12_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_19_io_mulInput = mac_11_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_19_io_addInput = mac_12_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_20_clock = clock;
  assign mac_12_20_reset = reset;
  assign mac_12_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_20_io_mulInput = mac_11_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_20_io_addInput = mac_12_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_21_clock = clock;
  assign mac_12_21_reset = reset;
  assign mac_12_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_21_io_mulInput = mac_11_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_21_io_addInput = mac_12_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_22_clock = clock;
  assign mac_12_22_reset = reset;
  assign mac_12_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_22_io_mulInput = mac_11_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_22_io_addInput = mac_12_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_23_clock = clock;
  assign mac_12_23_reset = reset;
  assign mac_12_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_23_io_mulInput = mac_11_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_23_io_addInput = mac_12_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_24_clock = clock;
  assign mac_12_24_reset = reset;
  assign mac_12_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_24_io_mulInput = mac_11_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_24_io_addInput = mac_12_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_25_clock = clock;
  assign mac_12_25_reset = reset;
  assign mac_12_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_25_io_mulInput = mac_11_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_25_io_addInput = mac_12_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_26_clock = clock;
  assign mac_12_26_reset = reset;
  assign mac_12_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_26_io_mulInput = mac_11_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_26_io_addInput = mac_12_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_27_clock = clock;
  assign mac_12_27_reset = reset;
  assign mac_12_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_27_io_mulInput = mac_11_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_27_io_addInput = mac_12_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_28_clock = clock;
  assign mac_12_28_reset = reset;
  assign mac_12_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_28_io_mulInput = mac_11_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_28_io_addInput = mac_12_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_29_clock = clock;
  assign mac_12_29_reset = reset;
  assign mac_12_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_29_io_mulInput = mac_11_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_29_io_addInput = mac_12_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_30_clock = clock;
  assign mac_12_30_reset = reset;
  assign mac_12_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_30_io_mulInput = mac_11_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_30_io_addInput = mac_12_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_12_31_clock = clock;
  assign mac_12_31_reset = reset;
  assign mac_12_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_12_31_io_mulInput = mac_11_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_12_31_io_addInput = mac_12_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_0_clock = clock;
  assign mac_13_0_reset = reset;
  assign mac_13_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_13_0_io_mulInput = mac_12_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_13_0_io_addInput = bias_13; // @[InnerSystolicArray.scala 57:27]
  assign mac_13_1_clock = clock;
  assign mac_13_1_reset = reset;
  assign mac_13_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_1_io_mulInput = mac_12_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_1_io_addInput = mac_13_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_2_clock = clock;
  assign mac_13_2_reset = reset;
  assign mac_13_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_2_io_mulInput = mac_12_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_2_io_addInput = mac_13_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_3_clock = clock;
  assign mac_13_3_reset = reset;
  assign mac_13_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_3_io_mulInput = mac_12_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_3_io_addInput = mac_13_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_4_clock = clock;
  assign mac_13_4_reset = reset;
  assign mac_13_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_4_io_mulInput = mac_12_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_4_io_addInput = mac_13_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_5_clock = clock;
  assign mac_13_5_reset = reset;
  assign mac_13_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_5_io_mulInput = mac_12_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_5_io_addInput = mac_13_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_6_clock = clock;
  assign mac_13_6_reset = reset;
  assign mac_13_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_6_io_mulInput = mac_12_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_6_io_addInput = mac_13_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_7_clock = clock;
  assign mac_13_7_reset = reset;
  assign mac_13_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_7_io_mulInput = mac_12_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_7_io_addInput = mac_13_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_8_clock = clock;
  assign mac_13_8_reset = reset;
  assign mac_13_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_8_io_mulInput = mac_12_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_8_io_addInput = mac_13_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_9_clock = clock;
  assign mac_13_9_reset = reset;
  assign mac_13_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_9_io_mulInput = mac_12_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_9_io_addInput = mac_13_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_10_clock = clock;
  assign mac_13_10_reset = reset;
  assign mac_13_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_10_io_mulInput = mac_12_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_10_io_addInput = mac_13_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_11_clock = clock;
  assign mac_13_11_reset = reset;
  assign mac_13_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_11_io_mulInput = mac_12_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_11_io_addInput = mac_13_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_12_clock = clock;
  assign mac_13_12_reset = reset;
  assign mac_13_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_12_io_mulInput = mac_12_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_12_io_addInput = mac_13_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_13_clock = clock;
  assign mac_13_13_reset = reset;
  assign mac_13_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_13_io_mulInput = mac_12_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_13_io_addInput = mac_13_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_14_clock = clock;
  assign mac_13_14_reset = reset;
  assign mac_13_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_14_io_mulInput = mac_12_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_14_io_addInput = mac_13_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_15_clock = clock;
  assign mac_13_15_reset = reset;
  assign mac_13_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_15_io_mulInput = mac_12_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_15_io_addInput = mac_13_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_16_clock = clock;
  assign mac_13_16_reset = reset;
  assign mac_13_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_16_io_mulInput = mac_12_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_16_io_addInput = mac_13_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_17_clock = clock;
  assign mac_13_17_reset = reset;
  assign mac_13_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_17_io_mulInput = mac_12_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_17_io_addInput = mac_13_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_18_clock = clock;
  assign mac_13_18_reset = reset;
  assign mac_13_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_18_io_mulInput = mac_12_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_18_io_addInput = mac_13_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_19_clock = clock;
  assign mac_13_19_reset = reset;
  assign mac_13_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_19_io_mulInput = mac_12_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_19_io_addInput = mac_13_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_20_clock = clock;
  assign mac_13_20_reset = reset;
  assign mac_13_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_20_io_mulInput = mac_12_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_20_io_addInput = mac_13_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_21_clock = clock;
  assign mac_13_21_reset = reset;
  assign mac_13_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_21_io_mulInput = mac_12_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_21_io_addInput = mac_13_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_22_clock = clock;
  assign mac_13_22_reset = reset;
  assign mac_13_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_22_io_mulInput = mac_12_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_22_io_addInput = mac_13_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_23_clock = clock;
  assign mac_13_23_reset = reset;
  assign mac_13_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_23_io_mulInput = mac_12_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_23_io_addInput = mac_13_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_24_clock = clock;
  assign mac_13_24_reset = reset;
  assign mac_13_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_24_io_mulInput = mac_12_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_24_io_addInput = mac_13_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_25_clock = clock;
  assign mac_13_25_reset = reset;
  assign mac_13_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_25_io_mulInput = mac_12_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_25_io_addInput = mac_13_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_26_clock = clock;
  assign mac_13_26_reset = reset;
  assign mac_13_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_26_io_mulInput = mac_12_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_26_io_addInput = mac_13_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_27_clock = clock;
  assign mac_13_27_reset = reset;
  assign mac_13_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_27_io_mulInput = mac_12_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_27_io_addInput = mac_13_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_28_clock = clock;
  assign mac_13_28_reset = reset;
  assign mac_13_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_28_io_mulInput = mac_12_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_28_io_addInput = mac_13_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_29_clock = clock;
  assign mac_13_29_reset = reset;
  assign mac_13_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_29_io_mulInput = mac_12_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_29_io_addInput = mac_13_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_30_clock = clock;
  assign mac_13_30_reset = reset;
  assign mac_13_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_30_io_mulInput = mac_12_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_30_io_addInput = mac_13_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_13_31_clock = clock;
  assign mac_13_31_reset = reset;
  assign mac_13_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_13_31_io_mulInput = mac_12_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_13_31_io_addInput = mac_13_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_0_clock = clock;
  assign mac_14_0_reset = reset;
  assign mac_14_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_14_0_io_mulInput = mac_13_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_14_0_io_addInput = bias_14; // @[InnerSystolicArray.scala 57:27]
  assign mac_14_1_clock = clock;
  assign mac_14_1_reset = reset;
  assign mac_14_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_1_io_mulInput = mac_13_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_1_io_addInput = mac_14_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_2_clock = clock;
  assign mac_14_2_reset = reset;
  assign mac_14_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_2_io_mulInput = mac_13_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_2_io_addInput = mac_14_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_3_clock = clock;
  assign mac_14_3_reset = reset;
  assign mac_14_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_3_io_mulInput = mac_13_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_3_io_addInput = mac_14_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_4_clock = clock;
  assign mac_14_4_reset = reset;
  assign mac_14_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_4_io_mulInput = mac_13_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_4_io_addInput = mac_14_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_5_clock = clock;
  assign mac_14_5_reset = reset;
  assign mac_14_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_5_io_mulInput = mac_13_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_5_io_addInput = mac_14_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_6_clock = clock;
  assign mac_14_6_reset = reset;
  assign mac_14_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_6_io_mulInput = mac_13_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_6_io_addInput = mac_14_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_7_clock = clock;
  assign mac_14_7_reset = reset;
  assign mac_14_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_7_io_mulInput = mac_13_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_7_io_addInput = mac_14_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_8_clock = clock;
  assign mac_14_8_reset = reset;
  assign mac_14_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_8_io_mulInput = mac_13_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_8_io_addInput = mac_14_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_9_clock = clock;
  assign mac_14_9_reset = reset;
  assign mac_14_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_9_io_mulInput = mac_13_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_9_io_addInput = mac_14_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_10_clock = clock;
  assign mac_14_10_reset = reset;
  assign mac_14_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_10_io_mulInput = mac_13_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_10_io_addInput = mac_14_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_11_clock = clock;
  assign mac_14_11_reset = reset;
  assign mac_14_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_11_io_mulInput = mac_13_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_11_io_addInput = mac_14_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_12_clock = clock;
  assign mac_14_12_reset = reset;
  assign mac_14_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_12_io_mulInput = mac_13_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_12_io_addInput = mac_14_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_13_clock = clock;
  assign mac_14_13_reset = reset;
  assign mac_14_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_13_io_mulInput = mac_13_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_13_io_addInput = mac_14_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_14_clock = clock;
  assign mac_14_14_reset = reset;
  assign mac_14_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_14_io_mulInput = mac_13_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_14_io_addInput = mac_14_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_15_clock = clock;
  assign mac_14_15_reset = reset;
  assign mac_14_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_15_io_mulInput = mac_13_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_15_io_addInput = mac_14_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_16_clock = clock;
  assign mac_14_16_reset = reset;
  assign mac_14_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_16_io_mulInput = mac_13_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_16_io_addInput = mac_14_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_17_clock = clock;
  assign mac_14_17_reset = reset;
  assign mac_14_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_17_io_mulInput = mac_13_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_17_io_addInput = mac_14_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_18_clock = clock;
  assign mac_14_18_reset = reset;
  assign mac_14_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_18_io_mulInput = mac_13_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_18_io_addInput = mac_14_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_19_clock = clock;
  assign mac_14_19_reset = reset;
  assign mac_14_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_19_io_mulInput = mac_13_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_19_io_addInput = mac_14_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_20_clock = clock;
  assign mac_14_20_reset = reset;
  assign mac_14_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_20_io_mulInput = mac_13_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_20_io_addInput = mac_14_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_21_clock = clock;
  assign mac_14_21_reset = reset;
  assign mac_14_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_21_io_mulInput = mac_13_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_21_io_addInput = mac_14_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_22_clock = clock;
  assign mac_14_22_reset = reset;
  assign mac_14_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_22_io_mulInput = mac_13_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_22_io_addInput = mac_14_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_23_clock = clock;
  assign mac_14_23_reset = reset;
  assign mac_14_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_23_io_mulInput = mac_13_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_23_io_addInput = mac_14_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_24_clock = clock;
  assign mac_14_24_reset = reset;
  assign mac_14_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_24_io_mulInput = mac_13_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_24_io_addInput = mac_14_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_25_clock = clock;
  assign mac_14_25_reset = reset;
  assign mac_14_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_25_io_mulInput = mac_13_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_25_io_addInput = mac_14_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_26_clock = clock;
  assign mac_14_26_reset = reset;
  assign mac_14_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_26_io_mulInput = mac_13_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_26_io_addInput = mac_14_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_27_clock = clock;
  assign mac_14_27_reset = reset;
  assign mac_14_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_27_io_mulInput = mac_13_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_27_io_addInput = mac_14_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_28_clock = clock;
  assign mac_14_28_reset = reset;
  assign mac_14_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_28_io_mulInput = mac_13_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_28_io_addInput = mac_14_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_29_clock = clock;
  assign mac_14_29_reset = reset;
  assign mac_14_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_29_io_mulInput = mac_13_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_29_io_addInput = mac_14_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_30_clock = clock;
  assign mac_14_30_reset = reset;
  assign mac_14_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_30_io_mulInput = mac_13_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_30_io_addInput = mac_14_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_14_31_clock = clock;
  assign mac_14_31_reset = reset;
  assign mac_14_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_14_31_io_mulInput = mac_13_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_14_31_io_addInput = mac_14_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_0_clock = clock;
  assign mac_15_0_reset = reset;
  assign mac_15_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_15_0_io_mulInput = mac_14_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_15_0_io_addInput = bias_15; // @[InnerSystolicArray.scala 57:27]
  assign mac_15_1_clock = clock;
  assign mac_15_1_reset = reset;
  assign mac_15_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_1_io_mulInput = mac_14_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_1_io_addInput = mac_15_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_2_clock = clock;
  assign mac_15_2_reset = reset;
  assign mac_15_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_2_io_mulInput = mac_14_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_2_io_addInput = mac_15_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_3_clock = clock;
  assign mac_15_3_reset = reset;
  assign mac_15_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_3_io_mulInput = mac_14_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_3_io_addInput = mac_15_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_4_clock = clock;
  assign mac_15_4_reset = reset;
  assign mac_15_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_4_io_mulInput = mac_14_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_4_io_addInput = mac_15_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_5_clock = clock;
  assign mac_15_5_reset = reset;
  assign mac_15_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_5_io_mulInput = mac_14_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_5_io_addInput = mac_15_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_6_clock = clock;
  assign mac_15_6_reset = reset;
  assign mac_15_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_6_io_mulInput = mac_14_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_6_io_addInput = mac_15_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_7_clock = clock;
  assign mac_15_7_reset = reset;
  assign mac_15_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_7_io_mulInput = mac_14_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_7_io_addInput = mac_15_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_8_clock = clock;
  assign mac_15_8_reset = reset;
  assign mac_15_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_8_io_mulInput = mac_14_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_8_io_addInput = mac_15_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_9_clock = clock;
  assign mac_15_9_reset = reset;
  assign mac_15_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_9_io_mulInput = mac_14_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_9_io_addInput = mac_15_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_10_clock = clock;
  assign mac_15_10_reset = reset;
  assign mac_15_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_10_io_mulInput = mac_14_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_10_io_addInput = mac_15_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_11_clock = clock;
  assign mac_15_11_reset = reset;
  assign mac_15_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_11_io_mulInput = mac_14_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_11_io_addInput = mac_15_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_12_clock = clock;
  assign mac_15_12_reset = reset;
  assign mac_15_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_12_io_mulInput = mac_14_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_12_io_addInput = mac_15_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_13_clock = clock;
  assign mac_15_13_reset = reset;
  assign mac_15_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_13_io_mulInput = mac_14_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_13_io_addInput = mac_15_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_14_clock = clock;
  assign mac_15_14_reset = reset;
  assign mac_15_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_14_io_mulInput = mac_14_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_14_io_addInput = mac_15_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_15_clock = clock;
  assign mac_15_15_reset = reset;
  assign mac_15_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_15_io_mulInput = mac_14_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_15_io_addInput = mac_15_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_16_clock = clock;
  assign mac_15_16_reset = reset;
  assign mac_15_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_16_io_mulInput = mac_14_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_16_io_addInput = mac_15_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_17_clock = clock;
  assign mac_15_17_reset = reset;
  assign mac_15_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_17_io_mulInput = mac_14_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_17_io_addInput = mac_15_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_18_clock = clock;
  assign mac_15_18_reset = reset;
  assign mac_15_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_18_io_mulInput = mac_14_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_18_io_addInput = mac_15_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_19_clock = clock;
  assign mac_15_19_reset = reset;
  assign mac_15_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_19_io_mulInput = mac_14_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_19_io_addInput = mac_15_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_20_clock = clock;
  assign mac_15_20_reset = reset;
  assign mac_15_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_20_io_mulInput = mac_14_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_20_io_addInput = mac_15_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_21_clock = clock;
  assign mac_15_21_reset = reset;
  assign mac_15_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_21_io_mulInput = mac_14_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_21_io_addInput = mac_15_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_22_clock = clock;
  assign mac_15_22_reset = reset;
  assign mac_15_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_22_io_mulInput = mac_14_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_22_io_addInput = mac_15_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_23_clock = clock;
  assign mac_15_23_reset = reset;
  assign mac_15_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_23_io_mulInput = mac_14_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_23_io_addInput = mac_15_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_24_clock = clock;
  assign mac_15_24_reset = reset;
  assign mac_15_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_24_io_mulInput = mac_14_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_24_io_addInput = mac_15_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_25_clock = clock;
  assign mac_15_25_reset = reset;
  assign mac_15_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_25_io_mulInput = mac_14_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_25_io_addInput = mac_15_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_26_clock = clock;
  assign mac_15_26_reset = reset;
  assign mac_15_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_26_io_mulInput = mac_14_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_26_io_addInput = mac_15_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_27_clock = clock;
  assign mac_15_27_reset = reset;
  assign mac_15_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_27_io_mulInput = mac_14_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_27_io_addInput = mac_15_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_28_clock = clock;
  assign mac_15_28_reset = reset;
  assign mac_15_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_28_io_mulInput = mac_14_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_28_io_addInput = mac_15_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_29_clock = clock;
  assign mac_15_29_reset = reset;
  assign mac_15_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_29_io_mulInput = mac_14_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_29_io_addInput = mac_15_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_30_clock = clock;
  assign mac_15_30_reset = reset;
  assign mac_15_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_30_io_mulInput = mac_14_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_30_io_addInput = mac_15_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_15_31_clock = clock;
  assign mac_15_31_reset = reset;
  assign mac_15_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_15_31_io_mulInput = mac_14_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_15_31_io_addInput = mac_15_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_0_clock = clock;
  assign mac_16_0_reset = reset;
  assign mac_16_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_16_0_io_mulInput = mac_15_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_16_0_io_addInput = bias_16; // @[InnerSystolicArray.scala 57:27]
  assign mac_16_1_clock = clock;
  assign mac_16_1_reset = reset;
  assign mac_16_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_1_io_mulInput = mac_15_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_1_io_addInput = mac_16_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_2_clock = clock;
  assign mac_16_2_reset = reset;
  assign mac_16_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_2_io_mulInput = mac_15_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_2_io_addInput = mac_16_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_3_clock = clock;
  assign mac_16_3_reset = reset;
  assign mac_16_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_3_io_mulInput = mac_15_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_3_io_addInput = mac_16_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_4_clock = clock;
  assign mac_16_4_reset = reset;
  assign mac_16_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_4_io_mulInput = mac_15_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_4_io_addInput = mac_16_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_5_clock = clock;
  assign mac_16_5_reset = reset;
  assign mac_16_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_5_io_mulInput = mac_15_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_5_io_addInput = mac_16_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_6_clock = clock;
  assign mac_16_6_reset = reset;
  assign mac_16_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_6_io_mulInput = mac_15_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_6_io_addInput = mac_16_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_7_clock = clock;
  assign mac_16_7_reset = reset;
  assign mac_16_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_7_io_mulInput = mac_15_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_7_io_addInput = mac_16_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_8_clock = clock;
  assign mac_16_8_reset = reset;
  assign mac_16_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_8_io_mulInput = mac_15_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_8_io_addInput = mac_16_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_9_clock = clock;
  assign mac_16_9_reset = reset;
  assign mac_16_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_9_io_mulInput = mac_15_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_9_io_addInput = mac_16_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_10_clock = clock;
  assign mac_16_10_reset = reset;
  assign mac_16_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_10_io_mulInput = mac_15_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_10_io_addInput = mac_16_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_11_clock = clock;
  assign mac_16_11_reset = reset;
  assign mac_16_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_11_io_mulInput = mac_15_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_11_io_addInput = mac_16_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_12_clock = clock;
  assign mac_16_12_reset = reset;
  assign mac_16_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_12_io_mulInput = mac_15_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_12_io_addInput = mac_16_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_13_clock = clock;
  assign mac_16_13_reset = reset;
  assign mac_16_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_13_io_mulInput = mac_15_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_13_io_addInput = mac_16_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_14_clock = clock;
  assign mac_16_14_reset = reset;
  assign mac_16_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_14_io_mulInput = mac_15_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_14_io_addInput = mac_16_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_15_clock = clock;
  assign mac_16_15_reset = reset;
  assign mac_16_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_15_io_mulInput = mac_15_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_15_io_addInput = mac_16_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_16_clock = clock;
  assign mac_16_16_reset = reset;
  assign mac_16_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_16_io_mulInput = mac_15_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_16_io_addInput = mac_16_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_17_clock = clock;
  assign mac_16_17_reset = reset;
  assign mac_16_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_17_io_mulInput = mac_15_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_17_io_addInput = mac_16_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_18_clock = clock;
  assign mac_16_18_reset = reset;
  assign mac_16_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_18_io_mulInput = mac_15_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_18_io_addInput = mac_16_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_19_clock = clock;
  assign mac_16_19_reset = reset;
  assign mac_16_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_19_io_mulInput = mac_15_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_19_io_addInput = mac_16_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_20_clock = clock;
  assign mac_16_20_reset = reset;
  assign mac_16_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_20_io_mulInput = mac_15_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_20_io_addInput = mac_16_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_21_clock = clock;
  assign mac_16_21_reset = reset;
  assign mac_16_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_21_io_mulInput = mac_15_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_21_io_addInput = mac_16_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_22_clock = clock;
  assign mac_16_22_reset = reset;
  assign mac_16_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_22_io_mulInput = mac_15_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_22_io_addInput = mac_16_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_23_clock = clock;
  assign mac_16_23_reset = reset;
  assign mac_16_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_23_io_mulInput = mac_15_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_23_io_addInput = mac_16_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_24_clock = clock;
  assign mac_16_24_reset = reset;
  assign mac_16_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_24_io_mulInput = mac_15_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_24_io_addInput = mac_16_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_25_clock = clock;
  assign mac_16_25_reset = reset;
  assign mac_16_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_25_io_mulInput = mac_15_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_25_io_addInput = mac_16_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_26_clock = clock;
  assign mac_16_26_reset = reset;
  assign mac_16_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_26_io_mulInput = mac_15_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_26_io_addInput = mac_16_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_27_clock = clock;
  assign mac_16_27_reset = reset;
  assign mac_16_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_27_io_mulInput = mac_15_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_27_io_addInput = mac_16_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_28_clock = clock;
  assign mac_16_28_reset = reset;
  assign mac_16_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_28_io_mulInput = mac_15_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_28_io_addInput = mac_16_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_29_clock = clock;
  assign mac_16_29_reset = reset;
  assign mac_16_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_29_io_mulInput = mac_15_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_29_io_addInput = mac_16_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_30_clock = clock;
  assign mac_16_30_reset = reset;
  assign mac_16_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_30_io_mulInput = mac_15_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_30_io_addInput = mac_16_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_16_31_clock = clock;
  assign mac_16_31_reset = reset;
  assign mac_16_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_16_31_io_mulInput = mac_15_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_16_31_io_addInput = mac_16_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_0_clock = clock;
  assign mac_17_0_reset = reset;
  assign mac_17_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_17_0_io_mulInput = mac_16_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_17_0_io_addInput = bias_17; // @[InnerSystolicArray.scala 57:27]
  assign mac_17_1_clock = clock;
  assign mac_17_1_reset = reset;
  assign mac_17_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_1_io_mulInput = mac_16_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_1_io_addInput = mac_17_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_2_clock = clock;
  assign mac_17_2_reset = reset;
  assign mac_17_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_2_io_mulInput = mac_16_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_2_io_addInput = mac_17_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_3_clock = clock;
  assign mac_17_3_reset = reset;
  assign mac_17_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_3_io_mulInput = mac_16_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_3_io_addInput = mac_17_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_4_clock = clock;
  assign mac_17_4_reset = reset;
  assign mac_17_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_4_io_mulInput = mac_16_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_4_io_addInput = mac_17_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_5_clock = clock;
  assign mac_17_5_reset = reset;
  assign mac_17_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_5_io_mulInput = mac_16_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_5_io_addInput = mac_17_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_6_clock = clock;
  assign mac_17_6_reset = reset;
  assign mac_17_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_6_io_mulInput = mac_16_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_6_io_addInput = mac_17_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_7_clock = clock;
  assign mac_17_7_reset = reset;
  assign mac_17_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_7_io_mulInput = mac_16_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_7_io_addInput = mac_17_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_8_clock = clock;
  assign mac_17_8_reset = reset;
  assign mac_17_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_8_io_mulInput = mac_16_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_8_io_addInput = mac_17_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_9_clock = clock;
  assign mac_17_9_reset = reset;
  assign mac_17_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_9_io_mulInput = mac_16_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_9_io_addInput = mac_17_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_10_clock = clock;
  assign mac_17_10_reset = reset;
  assign mac_17_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_10_io_mulInput = mac_16_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_10_io_addInput = mac_17_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_11_clock = clock;
  assign mac_17_11_reset = reset;
  assign mac_17_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_11_io_mulInput = mac_16_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_11_io_addInput = mac_17_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_12_clock = clock;
  assign mac_17_12_reset = reset;
  assign mac_17_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_12_io_mulInput = mac_16_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_12_io_addInput = mac_17_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_13_clock = clock;
  assign mac_17_13_reset = reset;
  assign mac_17_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_13_io_mulInput = mac_16_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_13_io_addInput = mac_17_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_14_clock = clock;
  assign mac_17_14_reset = reset;
  assign mac_17_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_14_io_mulInput = mac_16_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_14_io_addInput = mac_17_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_15_clock = clock;
  assign mac_17_15_reset = reset;
  assign mac_17_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_15_io_mulInput = mac_16_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_15_io_addInput = mac_17_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_16_clock = clock;
  assign mac_17_16_reset = reset;
  assign mac_17_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_16_io_mulInput = mac_16_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_16_io_addInput = mac_17_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_17_clock = clock;
  assign mac_17_17_reset = reset;
  assign mac_17_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_17_io_mulInput = mac_16_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_17_io_addInput = mac_17_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_18_clock = clock;
  assign mac_17_18_reset = reset;
  assign mac_17_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_18_io_mulInput = mac_16_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_18_io_addInput = mac_17_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_19_clock = clock;
  assign mac_17_19_reset = reset;
  assign mac_17_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_19_io_mulInput = mac_16_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_19_io_addInput = mac_17_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_20_clock = clock;
  assign mac_17_20_reset = reset;
  assign mac_17_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_20_io_mulInput = mac_16_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_20_io_addInput = mac_17_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_21_clock = clock;
  assign mac_17_21_reset = reset;
  assign mac_17_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_21_io_mulInput = mac_16_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_21_io_addInput = mac_17_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_22_clock = clock;
  assign mac_17_22_reset = reset;
  assign mac_17_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_22_io_mulInput = mac_16_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_22_io_addInput = mac_17_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_23_clock = clock;
  assign mac_17_23_reset = reset;
  assign mac_17_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_23_io_mulInput = mac_16_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_23_io_addInput = mac_17_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_24_clock = clock;
  assign mac_17_24_reset = reset;
  assign mac_17_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_24_io_mulInput = mac_16_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_24_io_addInput = mac_17_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_25_clock = clock;
  assign mac_17_25_reset = reset;
  assign mac_17_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_25_io_mulInput = mac_16_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_25_io_addInput = mac_17_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_26_clock = clock;
  assign mac_17_26_reset = reset;
  assign mac_17_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_26_io_mulInput = mac_16_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_26_io_addInput = mac_17_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_27_clock = clock;
  assign mac_17_27_reset = reset;
  assign mac_17_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_27_io_mulInput = mac_16_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_27_io_addInput = mac_17_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_28_clock = clock;
  assign mac_17_28_reset = reset;
  assign mac_17_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_28_io_mulInput = mac_16_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_28_io_addInput = mac_17_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_29_clock = clock;
  assign mac_17_29_reset = reset;
  assign mac_17_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_29_io_mulInput = mac_16_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_29_io_addInput = mac_17_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_30_clock = clock;
  assign mac_17_30_reset = reset;
  assign mac_17_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_30_io_mulInput = mac_16_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_30_io_addInput = mac_17_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_17_31_clock = clock;
  assign mac_17_31_reset = reset;
  assign mac_17_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_17_31_io_mulInput = mac_16_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_17_31_io_addInput = mac_17_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_0_clock = clock;
  assign mac_18_0_reset = reset;
  assign mac_18_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_18_0_io_mulInput = mac_17_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_18_0_io_addInput = bias_18; // @[InnerSystolicArray.scala 57:27]
  assign mac_18_1_clock = clock;
  assign mac_18_1_reset = reset;
  assign mac_18_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_1_io_mulInput = mac_17_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_1_io_addInput = mac_18_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_2_clock = clock;
  assign mac_18_2_reset = reset;
  assign mac_18_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_2_io_mulInput = mac_17_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_2_io_addInput = mac_18_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_3_clock = clock;
  assign mac_18_3_reset = reset;
  assign mac_18_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_3_io_mulInput = mac_17_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_3_io_addInput = mac_18_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_4_clock = clock;
  assign mac_18_4_reset = reset;
  assign mac_18_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_4_io_mulInput = mac_17_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_4_io_addInput = mac_18_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_5_clock = clock;
  assign mac_18_5_reset = reset;
  assign mac_18_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_5_io_mulInput = mac_17_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_5_io_addInput = mac_18_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_6_clock = clock;
  assign mac_18_6_reset = reset;
  assign mac_18_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_6_io_mulInput = mac_17_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_6_io_addInput = mac_18_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_7_clock = clock;
  assign mac_18_7_reset = reset;
  assign mac_18_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_7_io_mulInput = mac_17_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_7_io_addInput = mac_18_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_8_clock = clock;
  assign mac_18_8_reset = reset;
  assign mac_18_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_8_io_mulInput = mac_17_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_8_io_addInput = mac_18_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_9_clock = clock;
  assign mac_18_9_reset = reset;
  assign mac_18_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_9_io_mulInput = mac_17_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_9_io_addInput = mac_18_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_10_clock = clock;
  assign mac_18_10_reset = reset;
  assign mac_18_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_10_io_mulInput = mac_17_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_10_io_addInput = mac_18_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_11_clock = clock;
  assign mac_18_11_reset = reset;
  assign mac_18_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_11_io_mulInput = mac_17_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_11_io_addInput = mac_18_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_12_clock = clock;
  assign mac_18_12_reset = reset;
  assign mac_18_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_12_io_mulInput = mac_17_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_12_io_addInput = mac_18_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_13_clock = clock;
  assign mac_18_13_reset = reset;
  assign mac_18_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_13_io_mulInput = mac_17_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_13_io_addInput = mac_18_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_14_clock = clock;
  assign mac_18_14_reset = reset;
  assign mac_18_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_14_io_mulInput = mac_17_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_14_io_addInput = mac_18_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_15_clock = clock;
  assign mac_18_15_reset = reset;
  assign mac_18_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_15_io_mulInput = mac_17_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_15_io_addInput = mac_18_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_16_clock = clock;
  assign mac_18_16_reset = reset;
  assign mac_18_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_16_io_mulInput = mac_17_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_16_io_addInput = mac_18_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_17_clock = clock;
  assign mac_18_17_reset = reset;
  assign mac_18_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_17_io_mulInput = mac_17_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_17_io_addInput = mac_18_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_18_clock = clock;
  assign mac_18_18_reset = reset;
  assign mac_18_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_18_io_mulInput = mac_17_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_18_io_addInput = mac_18_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_19_clock = clock;
  assign mac_18_19_reset = reset;
  assign mac_18_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_19_io_mulInput = mac_17_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_19_io_addInput = mac_18_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_20_clock = clock;
  assign mac_18_20_reset = reset;
  assign mac_18_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_20_io_mulInput = mac_17_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_20_io_addInput = mac_18_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_21_clock = clock;
  assign mac_18_21_reset = reset;
  assign mac_18_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_21_io_mulInput = mac_17_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_21_io_addInput = mac_18_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_22_clock = clock;
  assign mac_18_22_reset = reset;
  assign mac_18_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_22_io_mulInput = mac_17_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_22_io_addInput = mac_18_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_23_clock = clock;
  assign mac_18_23_reset = reset;
  assign mac_18_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_23_io_mulInput = mac_17_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_23_io_addInput = mac_18_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_24_clock = clock;
  assign mac_18_24_reset = reset;
  assign mac_18_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_24_io_mulInput = mac_17_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_24_io_addInput = mac_18_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_25_clock = clock;
  assign mac_18_25_reset = reset;
  assign mac_18_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_25_io_mulInput = mac_17_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_25_io_addInput = mac_18_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_26_clock = clock;
  assign mac_18_26_reset = reset;
  assign mac_18_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_26_io_mulInput = mac_17_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_26_io_addInput = mac_18_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_27_clock = clock;
  assign mac_18_27_reset = reset;
  assign mac_18_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_27_io_mulInput = mac_17_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_27_io_addInput = mac_18_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_28_clock = clock;
  assign mac_18_28_reset = reset;
  assign mac_18_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_28_io_mulInput = mac_17_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_28_io_addInput = mac_18_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_29_clock = clock;
  assign mac_18_29_reset = reset;
  assign mac_18_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_29_io_mulInput = mac_17_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_29_io_addInput = mac_18_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_30_clock = clock;
  assign mac_18_30_reset = reset;
  assign mac_18_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_30_io_mulInput = mac_17_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_30_io_addInput = mac_18_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_18_31_clock = clock;
  assign mac_18_31_reset = reset;
  assign mac_18_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_18_31_io_mulInput = mac_17_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_18_31_io_addInput = mac_18_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_0_clock = clock;
  assign mac_19_0_reset = reset;
  assign mac_19_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_19_0_io_mulInput = mac_18_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_19_0_io_addInput = bias_19; // @[InnerSystolicArray.scala 57:27]
  assign mac_19_1_clock = clock;
  assign mac_19_1_reset = reset;
  assign mac_19_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_1_io_mulInput = mac_18_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_1_io_addInput = mac_19_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_2_clock = clock;
  assign mac_19_2_reset = reset;
  assign mac_19_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_2_io_mulInput = mac_18_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_2_io_addInput = mac_19_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_3_clock = clock;
  assign mac_19_3_reset = reset;
  assign mac_19_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_3_io_mulInput = mac_18_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_3_io_addInput = mac_19_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_4_clock = clock;
  assign mac_19_4_reset = reset;
  assign mac_19_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_4_io_mulInput = mac_18_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_4_io_addInput = mac_19_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_5_clock = clock;
  assign mac_19_5_reset = reset;
  assign mac_19_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_5_io_mulInput = mac_18_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_5_io_addInput = mac_19_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_6_clock = clock;
  assign mac_19_6_reset = reset;
  assign mac_19_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_6_io_mulInput = mac_18_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_6_io_addInput = mac_19_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_7_clock = clock;
  assign mac_19_7_reset = reset;
  assign mac_19_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_7_io_mulInput = mac_18_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_7_io_addInput = mac_19_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_8_clock = clock;
  assign mac_19_8_reset = reset;
  assign mac_19_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_8_io_mulInput = mac_18_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_8_io_addInput = mac_19_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_9_clock = clock;
  assign mac_19_9_reset = reset;
  assign mac_19_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_9_io_mulInput = mac_18_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_9_io_addInput = mac_19_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_10_clock = clock;
  assign mac_19_10_reset = reset;
  assign mac_19_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_10_io_mulInput = mac_18_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_10_io_addInput = mac_19_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_11_clock = clock;
  assign mac_19_11_reset = reset;
  assign mac_19_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_11_io_mulInput = mac_18_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_11_io_addInput = mac_19_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_12_clock = clock;
  assign mac_19_12_reset = reset;
  assign mac_19_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_12_io_mulInput = mac_18_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_12_io_addInput = mac_19_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_13_clock = clock;
  assign mac_19_13_reset = reset;
  assign mac_19_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_13_io_mulInput = mac_18_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_13_io_addInput = mac_19_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_14_clock = clock;
  assign mac_19_14_reset = reset;
  assign mac_19_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_14_io_mulInput = mac_18_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_14_io_addInput = mac_19_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_15_clock = clock;
  assign mac_19_15_reset = reset;
  assign mac_19_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_15_io_mulInput = mac_18_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_15_io_addInput = mac_19_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_16_clock = clock;
  assign mac_19_16_reset = reset;
  assign mac_19_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_16_io_mulInput = mac_18_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_16_io_addInput = mac_19_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_17_clock = clock;
  assign mac_19_17_reset = reset;
  assign mac_19_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_17_io_mulInput = mac_18_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_17_io_addInput = mac_19_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_18_clock = clock;
  assign mac_19_18_reset = reset;
  assign mac_19_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_18_io_mulInput = mac_18_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_18_io_addInput = mac_19_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_19_clock = clock;
  assign mac_19_19_reset = reset;
  assign mac_19_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_19_io_mulInput = mac_18_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_19_io_addInput = mac_19_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_20_clock = clock;
  assign mac_19_20_reset = reset;
  assign mac_19_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_20_io_mulInput = mac_18_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_20_io_addInput = mac_19_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_21_clock = clock;
  assign mac_19_21_reset = reset;
  assign mac_19_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_21_io_mulInput = mac_18_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_21_io_addInput = mac_19_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_22_clock = clock;
  assign mac_19_22_reset = reset;
  assign mac_19_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_22_io_mulInput = mac_18_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_22_io_addInput = mac_19_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_23_clock = clock;
  assign mac_19_23_reset = reset;
  assign mac_19_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_23_io_mulInput = mac_18_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_23_io_addInput = mac_19_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_24_clock = clock;
  assign mac_19_24_reset = reset;
  assign mac_19_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_24_io_mulInput = mac_18_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_24_io_addInput = mac_19_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_25_clock = clock;
  assign mac_19_25_reset = reset;
  assign mac_19_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_25_io_mulInput = mac_18_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_25_io_addInput = mac_19_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_26_clock = clock;
  assign mac_19_26_reset = reset;
  assign mac_19_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_26_io_mulInput = mac_18_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_26_io_addInput = mac_19_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_27_clock = clock;
  assign mac_19_27_reset = reset;
  assign mac_19_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_27_io_mulInput = mac_18_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_27_io_addInput = mac_19_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_28_clock = clock;
  assign mac_19_28_reset = reset;
  assign mac_19_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_28_io_mulInput = mac_18_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_28_io_addInput = mac_19_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_29_clock = clock;
  assign mac_19_29_reset = reset;
  assign mac_19_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_29_io_mulInput = mac_18_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_29_io_addInput = mac_19_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_30_clock = clock;
  assign mac_19_30_reset = reset;
  assign mac_19_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_30_io_mulInput = mac_18_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_30_io_addInput = mac_19_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_19_31_clock = clock;
  assign mac_19_31_reset = reset;
  assign mac_19_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_19_31_io_mulInput = mac_18_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_19_31_io_addInput = mac_19_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_0_clock = clock;
  assign mac_20_0_reset = reset;
  assign mac_20_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_20_0_io_mulInput = mac_19_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_20_0_io_addInput = bias_20; // @[InnerSystolicArray.scala 57:27]
  assign mac_20_1_clock = clock;
  assign mac_20_1_reset = reset;
  assign mac_20_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_1_io_mulInput = mac_19_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_1_io_addInput = mac_20_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_2_clock = clock;
  assign mac_20_2_reset = reset;
  assign mac_20_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_2_io_mulInput = mac_19_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_2_io_addInput = mac_20_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_3_clock = clock;
  assign mac_20_3_reset = reset;
  assign mac_20_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_3_io_mulInput = mac_19_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_3_io_addInput = mac_20_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_4_clock = clock;
  assign mac_20_4_reset = reset;
  assign mac_20_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_4_io_mulInput = mac_19_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_4_io_addInput = mac_20_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_5_clock = clock;
  assign mac_20_5_reset = reset;
  assign mac_20_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_5_io_mulInput = mac_19_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_5_io_addInput = mac_20_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_6_clock = clock;
  assign mac_20_6_reset = reset;
  assign mac_20_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_6_io_mulInput = mac_19_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_6_io_addInput = mac_20_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_7_clock = clock;
  assign mac_20_7_reset = reset;
  assign mac_20_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_7_io_mulInput = mac_19_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_7_io_addInput = mac_20_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_8_clock = clock;
  assign mac_20_8_reset = reset;
  assign mac_20_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_8_io_mulInput = mac_19_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_8_io_addInput = mac_20_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_9_clock = clock;
  assign mac_20_9_reset = reset;
  assign mac_20_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_9_io_mulInput = mac_19_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_9_io_addInput = mac_20_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_10_clock = clock;
  assign mac_20_10_reset = reset;
  assign mac_20_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_10_io_mulInput = mac_19_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_10_io_addInput = mac_20_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_11_clock = clock;
  assign mac_20_11_reset = reset;
  assign mac_20_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_11_io_mulInput = mac_19_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_11_io_addInput = mac_20_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_12_clock = clock;
  assign mac_20_12_reset = reset;
  assign mac_20_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_12_io_mulInput = mac_19_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_12_io_addInput = mac_20_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_13_clock = clock;
  assign mac_20_13_reset = reset;
  assign mac_20_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_13_io_mulInput = mac_19_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_13_io_addInput = mac_20_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_14_clock = clock;
  assign mac_20_14_reset = reset;
  assign mac_20_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_14_io_mulInput = mac_19_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_14_io_addInput = mac_20_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_15_clock = clock;
  assign mac_20_15_reset = reset;
  assign mac_20_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_15_io_mulInput = mac_19_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_15_io_addInput = mac_20_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_16_clock = clock;
  assign mac_20_16_reset = reset;
  assign mac_20_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_16_io_mulInput = mac_19_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_16_io_addInput = mac_20_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_17_clock = clock;
  assign mac_20_17_reset = reset;
  assign mac_20_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_17_io_mulInput = mac_19_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_17_io_addInput = mac_20_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_18_clock = clock;
  assign mac_20_18_reset = reset;
  assign mac_20_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_18_io_mulInput = mac_19_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_18_io_addInput = mac_20_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_19_clock = clock;
  assign mac_20_19_reset = reset;
  assign mac_20_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_19_io_mulInput = mac_19_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_19_io_addInput = mac_20_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_20_clock = clock;
  assign mac_20_20_reset = reset;
  assign mac_20_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_20_io_mulInput = mac_19_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_20_io_addInput = mac_20_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_21_clock = clock;
  assign mac_20_21_reset = reset;
  assign mac_20_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_21_io_mulInput = mac_19_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_21_io_addInput = mac_20_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_22_clock = clock;
  assign mac_20_22_reset = reset;
  assign mac_20_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_22_io_mulInput = mac_19_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_22_io_addInput = mac_20_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_23_clock = clock;
  assign mac_20_23_reset = reset;
  assign mac_20_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_23_io_mulInput = mac_19_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_23_io_addInput = mac_20_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_24_clock = clock;
  assign mac_20_24_reset = reset;
  assign mac_20_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_24_io_mulInput = mac_19_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_24_io_addInput = mac_20_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_25_clock = clock;
  assign mac_20_25_reset = reset;
  assign mac_20_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_25_io_mulInput = mac_19_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_25_io_addInput = mac_20_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_26_clock = clock;
  assign mac_20_26_reset = reset;
  assign mac_20_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_26_io_mulInput = mac_19_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_26_io_addInput = mac_20_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_27_clock = clock;
  assign mac_20_27_reset = reset;
  assign mac_20_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_27_io_mulInput = mac_19_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_27_io_addInput = mac_20_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_28_clock = clock;
  assign mac_20_28_reset = reset;
  assign mac_20_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_28_io_mulInput = mac_19_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_28_io_addInput = mac_20_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_29_clock = clock;
  assign mac_20_29_reset = reset;
  assign mac_20_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_29_io_mulInput = mac_19_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_29_io_addInput = mac_20_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_30_clock = clock;
  assign mac_20_30_reset = reset;
  assign mac_20_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_30_io_mulInput = mac_19_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_30_io_addInput = mac_20_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_20_31_clock = clock;
  assign mac_20_31_reset = reset;
  assign mac_20_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_20_31_io_mulInput = mac_19_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_20_31_io_addInput = mac_20_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_0_clock = clock;
  assign mac_21_0_reset = reset;
  assign mac_21_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_21_0_io_mulInput = mac_20_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_21_0_io_addInput = bias_21; // @[InnerSystolicArray.scala 57:27]
  assign mac_21_1_clock = clock;
  assign mac_21_1_reset = reset;
  assign mac_21_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_1_io_mulInput = mac_20_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_1_io_addInput = mac_21_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_2_clock = clock;
  assign mac_21_2_reset = reset;
  assign mac_21_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_2_io_mulInput = mac_20_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_2_io_addInput = mac_21_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_3_clock = clock;
  assign mac_21_3_reset = reset;
  assign mac_21_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_3_io_mulInput = mac_20_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_3_io_addInput = mac_21_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_4_clock = clock;
  assign mac_21_4_reset = reset;
  assign mac_21_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_4_io_mulInput = mac_20_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_4_io_addInput = mac_21_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_5_clock = clock;
  assign mac_21_5_reset = reset;
  assign mac_21_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_5_io_mulInput = mac_20_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_5_io_addInput = mac_21_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_6_clock = clock;
  assign mac_21_6_reset = reset;
  assign mac_21_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_6_io_mulInput = mac_20_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_6_io_addInput = mac_21_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_7_clock = clock;
  assign mac_21_7_reset = reset;
  assign mac_21_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_7_io_mulInput = mac_20_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_7_io_addInput = mac_21_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_8_clock = clock;
  assign mac_21_8_reset = reset;
  assign mac_21_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_8_io_mulInput = mac_20_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_8_io_addInput = mac_21_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_9_clock = clock;
  assign mac_21_9_reset = reset;
  assign mac_21_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_9_io_mulInput = mac_20_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_9_io_addInput = mac_21_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_10_clock = clock;
  assign mac_21_10_reset = reset;
  assign mac_21_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_10_io_mulInput = mac_20_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_10_io_addInput = mac_21_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_11_clock = clock;
  assign mac_21_11_reset = reset;
  assign mac_21_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_11_io_mulInput = mac_20_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_11_io_addInput = mac_21_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_12_clock = clock;
  assign mac_21_12_reset = reset;
  assign mac_21_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_12_io_mulInput = mac_20_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_12_io_addInput = mac_21_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_13_clock = clock;
  assign mac_21_13_reset = reset;
  assign mac_21_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_13_io_mulInput = mac_20_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_13_io_addInput = mac_21_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_14_clock = clock;
  assign mac_21_14_reset = reset;
  assign mac_21_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_14_io_mulInput = mac_20_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_14_io_addInput = mac_21_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_15_clock = clock;
  assign mac_21_15_reset = reset;
  assign mac_21_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_15_io_mulInput = mac_20_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_15_io_addInput = mac_21_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_16_clock = clock;
  assign mac_21_16_reset = reset;
  assign mac_21_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_16_io_mulInput = mac_20_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_16_io_addInput = mac_21_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_17_clock = clock;
  assign mac_21_17_reset = reset;
  assign mac_21_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_17_io_mulInput = mac_20_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_17_io_addInput = mac_21_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_18_clock = clock;
  assign mac_21_18_reset = reset;
  assign mac_21_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_18_io_mulInput = mac_20_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_18_io_addInput = mac_21_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_19_clock = clock;
  assign mac_21_19_reset = reset;
  assign mac_21_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_19_io_mulInput = mac_20_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_19_io_addInput = mac_21_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_20_clock = clock;
  assign mac_21_20_reset = reset;
  assign mac_21_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_20_io_mulInput = mac_20_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_20_io_addInput = mac_21_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_21_clock = clock;
  assign mac_21_21_reset = reset;
  assign mac_21_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_21_io_mulInput = mac_20_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_21_io_addInput = mac_21_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_22_clock = clock;
  assign mac_21_22_reset = reset;
  assign mac_21_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_22_io_mulInput = mac_20_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_22_io_addInput = mac_21_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_23_clock = clock;
  assign mac_21_23_reset = reset;
  assign mac_21_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_23_io_mulInput = mac_20_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_23_io_addInput = mac_21_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_24_clock = clock;
  assign mac_21_24_reset = reset;
  assign mac_21_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_24_io_mulInput = mac_20_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_24_io_addInput = mac_21_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_25_clock = clock;
  assign mac_21_25_reset = reset;
  assign mac_21_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_25_io_mulInput = mac_20_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_25_io_addInput = mac_21_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_26_clock = clock;
  assign mac_21_26_reset = reset;
  assign mac_21_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_26_io_mulInput = mac_20_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_26_io_addInput = mac_21_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_27_clock = clock;
  assign mac_21_27_reset = reset;
  assign mac_21_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_27_io_mulInput = mac_20_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_27_io_addInput = mac_21_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_28_clock = clock;
  assign mac_21_28_reset = reset;
  assign mac_21_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_28_io_mulInput = mac_20_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_28_io_addInput = mac_21_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_29_clock = clock;
  assign mac_21_29_reset = reset;
  assign mac_21_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_29_io_mulInput = mac_20_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_29_io_addInput = mac_21_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_30_clock = clock;
  assign mac_21_30_reset = reset;
  assign mac_21_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_30_io_mulInput = mac_20_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_30_io_addInput = mac_21_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_21_31_clock = clock;
  assign mac_21_31_reset = reset;
  assign mac_21_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_21_31_io_mulInput = mac_20_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_21_31_io_addInput = mac_21_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_0_clock = clock;
  assign mac_22_0_reset = reset;
  assign mac_22_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_22_0_io_mulInput = mac_21_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_22_0_io_addInput = bias_22; // @[InnerSystolicArray.scala 57:27]
  assign mac_22_1_clock = clock;
  assign mac_22_1_reset = reset;
  assign mac_22_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_1_io_mulInput = mac_21_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_1_io_addInput = mac_22_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_2_clock = clock;
  assign mac_22_2_reset = reset;
  assign mac_22_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_2_io_mulInput = mac_21_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_2_io_addInput = mac_22_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_3_clock = clock;
  assign mac_22_3_reset = reset;
  assign mac_22_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_3_io_mulInput = mac_21_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_3_io_addInput = mac_22_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_4_clock = clock;
  assign mac_22_4_reset = reset;
  assign mac_22_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_4_io_mulInput = mac_21_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_4_io_addInput = mac_22_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_5_clock = clock;
  assign mac_22_5_reset = reset;
  assign mac_22_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_5_io_mulInput = mac_21_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_5_io_addInput = mac_22_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_6_clock = clock;
  assign mac_22_6_reset = reset;
  assign mac_22_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_6_io_mulInput = mac_21_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_6_io_addInput = mac_22_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_7_clock = clock;
  assign mac_22_7_reset = reset;
  assign mac_22_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_7_io_mulInput = mac_21_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_7_io_addInput = mac_22_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_8_clock = clock;
  assign mac_22_8_reset = reset;
  assign mac_22_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_8_io_mulInput = mac_21_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_8_io_addInput = mac_22_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_9_clock = clock;
  assign mac_22_9_reset = reset;
  assign mac_22_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_9_io_mulInput = mac_21_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_9_io_addInput = mac_22_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_10_clock = clock;
  assign mac_22_10_reset = reset;
  assign mac_22_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_10_io_mulInput = mac_21_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_10_io_addInput = mac_22_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_11_clock = clock;
  assign mac_22_11_reset = reset;
  assign mac_22_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_11_io_mulInput = mac_21_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_11_io_addInput = mac_22_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_12_clock = clock;
  assign mac_22_12_reset = reset;
  assign mac_22_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_12_io_mulInput = mac_21_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_12_io_addInput = mac_22_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_13_clock = clock;
  assign mac_22_13_reset = reset;
  assign mac_22_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_13_io_mulInput = mac_21_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_13_io_addInput = mac_22_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_14_clock = clock;
  assign mac_22_14_reset = reset;
  assign mac_22_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_14_io_mulInput = mac_21_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_14_io_addInput = mac_22_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_15_clock = clock;
  assign mac_22_15_reset = reset;
  assign mac_22_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_15_io_mulInput = mac_21_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_15_io_addInput = mac_22_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_16_clock = clock;
  assign mac_22_16_reset = reset;
  assign mac_22_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_16_io_mulInput = mac_21_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_16_io_addInput = mac_22_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_17_clock = clock;
  assign mac_22_17_reset = reset;
  assign mac_22_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_17_io_mulInput = mac_21_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_17_io_addInput = mac_22_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_18_clock = clock;
  assign mac_22_18_reset = reset;
  assign mac_22_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_18_io_mulInput = mac_21_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_18_io_addInput = mac_22_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_19_clock = clock;
  assign mac_22_19_reset = reset;
  assign mac_22_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_19_io_mulInput = mac_21_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_19_io_addInput = mac_22_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_20_clock = clock;
  assign mac_22_20_reset = reset;
  assign mac_22_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_20_io_mulInput = mac_21_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_20_io_addInput = mac_22_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_21_clock = clock;
  assign mac_22_21_reset = reset;
  assign mac_22_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_21_io_mulInput = mac_21_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_21_io_addInput = mac_22_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_22_clock = clock;
  assign mac_22_22_reset = reset;
  assign mac_22_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_22_io_mulInput = mac_21_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_22_io_addInput = mac_22_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_23_clock = clock;
  assign mac_22_23_reset = reset;
  assign mac_22_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_23_io_mulInput = mac_21_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_23_io_addInput = mac_22_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_24_clock = clock;
  assign mac_22_24_reset = reset;
  assign mac_22_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_24_io_mulInput = mac_21_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_24_io_addInput = mac_22_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_25_clock = clock;
  assign mac_22_25_reset = reset;
  assign mac_22_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_25_io_mulInput = mac_21_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_25_io_addInput = mac_22_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_26_clock = clock;
  assign mac_22_26_reset = reset;
  assign mac_22_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_26_io_mulInput = mac_21_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_26_io_addInput = mac_22_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_27_clock = clock;
  assign mac_22_27_reset = reset;
  assign mac_22_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_27_io_mulInput = mac_21_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_27_io_addInput = mac_22_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_28_clock = clock;
  assign mac_22_28_reset = reset;
  assign mac_22_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_28_io_mulInput = mac_21_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_28_io_addInput = mac_22_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_29_clock = clock;
  assign mac_22_29_reset = reset;
  assign mac_22_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_29_io_mulInput = mac_21_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_29_io_addInput = mac_22_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_30_clock = clock;
  assign mac_22_30_reset = reset;
  assign mac_22_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_30_io_mulInput = mac_21_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_30_io_addInput = mac_22_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_22_31_clock = clock;
  assign mac_22_31_reset = reset;
  assign mac_22_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_22_31_io_mulInput = mac_21_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_22_31_io_addInput = mac_22_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_0_clock = clock;
  assign mac_23_0_reset = reset;
  assign mac_23_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_23_0_io_mulInput = mac_22_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_23_0_io_addInput = bias_23; // @[InnerSystolicArray.scala 57:27]
  assign mac_23_1_clock = clock;
  assign mac_23_1_reset = reset;
  assign mac_23_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_1_io_mulInput = mac_22_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_1_io_addInput = mac_23_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_2_clock = clock;
  assign mac_23_2_reset = reset;
  assign mac_23_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_2_io_mulInput = mac_22_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_2_io_addInput = mac_23_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_3_clock = clock;
  assign mac_23_3_reset = reset;
  assign mac_23_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_3_io_mulInput = mac_22_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_3_io_addInput = mac_23_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_4_clock = clock;
  assign mac_23_4_reset = reset;
  assign mac_23_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_4_io_mulInput = mac_22_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_4_io_addInput = mac_23_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_5_clock = clock;
  assign mac_23_5_reset = reset;
  assign mac_23_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_5_io_mulInput = mac_22_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_5_io_addInput = mac_23_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_6_clock = clock;
  assign mac_23_6_reset = reset;
  assign mac_23_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_6_io_mulInput = mac_22_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_6_io_addInput = mac_23_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_7_clock = clock;
  assign mac_23_7_reset = reset;
  assign mac_23_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_7_io_mulInput = mac_22_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_7_io_addInput = mac_23_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_8_clock = clock;
  assign mac_23_8_reset = reset;
  assign mac_23_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_8_io_mulInput = mac_22_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_8_io_addInput = mac_23_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_9_clock = clock;
  assign mac_23_9_reset = reset;
  assign mac_23_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_9_io_mulInput = mac_22_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_9_io_addInput = mac_23_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_10_clock = clock;
  assign mac_23_10_reset = reset;
  assign mac_23_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_10_io_mulInput = mac_22_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_10_io_addInput = mac_23_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_11_clock = clock;
  assign mac_23_11_reset = reset;
  assign mac_23_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_11_io_mulInput = mac_22_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_11_io_addInput = mac_23_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_12_clock = clock;
  assign mac_23_12_reset = reset;
  assign mac_23_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_12_io_mulInput = mac_22_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_12_io_addInput = mac_23_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_13_clock = clock;
  assign mac_23_13_reset = reset;
  assign mac_23_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_13_io_mulInput = mac_22_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_13_io_addInput = mac_23_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_14_clock = clock;
  assign mac_23_14_reset = reset;
  assign mac_23_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_14_io_mulInput = mac_22_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_14_io_addInput = mac_23_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_15_clock = clock;
  assign mac_23_15_reset = reset;
  assign mac_23_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_15_io_mulInput = mac_22_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_15_io_addInput = mac_23_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_16_clock = clock;
  assign mac_23_16_reset = reset;
  assign mac_23_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_16_io_mulInput = mac_22_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_16_io_addInput = mac_23_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_17_clock = clock;
  assign mac_23_17_reset = reset;
  assign mac_23_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_17_io_mulInput = mac_22_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_17_io_addInput = mac_23_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_18_clock = clock;
  assign mac_23_18_reset = reset;
  assign mac_23_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_18_io_mulInput = mac_22_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_18_io_addInput = mac_23_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_19_clock = clock;
  assign mac_23_19_reset = reset;
  assign mac_23_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_19_io_mulInput = mac_22_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_19_io_addInput = mac_23_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_20_clock = clock;
  assign mac_23_20_reset = reset;
  assign mac_23_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_20_io_mulInput = mac_22_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_20_io_addInput = mac_23_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_21_clock = clock;
  assign mac_23_21_reset = reset;
  assign mac_23_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_21_io_mulInput = mac_22_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_21_io_addInput = mac_23_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_22_clock = clock;
  assign mac_23_22_reset = reset;
  assign mac_23_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_22_io_mulInput = mac_22_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_22_io_addInput = mac_23_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_23_clock = clock;
  assign mac_23_23_reset = reset;
  assign mac_23_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_23_io_mulInput = mac_22_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_23_io_addInput = mac_23_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_24_clock = clock;
  assign mac_23_24_reset = reset;
  assign mac_23_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_24_io_mulInput = mac_22_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_24_io_addInput = mac_23_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_25_clock = clock;
  assign mac_23_25_reset = reset;
  assign mac_23_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_25_io_mulInput = mac_22_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_25_io_addInput = mac_23_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_26_clock = clock;
  assign mac_23_26_reset = reset;
  assign mac_23_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_26_io_mulInput = mac_22_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_26_io_addInput = mac_23_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_27_clock = clock;
  assign mac_23_27_reset = reset;
  assign mac_23_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_27_io_mulInput = mac_22_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_27_io_addInput = mac_23_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_28_clock = clock;
  assign mac_23_28_reset = reset;
  assign mac_23_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_28_io_mulInput = mac_22_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_28_io_addInput = mac_23_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_29_clock = clock;
  assign mac_23_29_reset = reset;
  assign mac_23_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_29_io_mulInput = mac_22_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_29_io_addInput = mac_23_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_30_clock = clock;
  assign mac_23_30_reset = reset;
  assign mac_23_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_30_io_mulInput = mac_22_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_30_io_addInput = mac_23_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_23_31_clock = clock;
  assign mac_23_31_reset = reset;
  assign mac_23_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_23_31_io_mulInput = mac_22_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_23_31_io_addInput = mac_23_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_0_clock = clock;
  assign mac_24_0_reset = reset;
  assign mac_24_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_24_0_io_mulInput = mac_23_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_24_0_io_addInput = bias_24; // @[InnerSystolicArray.scala 57:27]
  assign mac_24_1_clock = clock;
  assign mac_24_1_reset = reset;
  assign mac_24_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_1_io_mulInput = mac_23_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_1_io_addInput = mac_24_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_2_clock = clock;
  assign mac_24_2_reset = reset;
  assign mac_24_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_2_io_mulInput = mac_23_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_2_io_addInput = mac_24_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_3_clock = clock;
  assign mac_24_3_reset = reset;
  assign mac_24_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_3_io_mulInput = mac_23_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_3_io_addInput = mac_24_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_4_clock = clock;
  assign mac_24_4_reset = reset;
  assign mac_24_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_4_io_mulInput = mac_23_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_4_io_addInput = mac_24_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_5_clock = clock;
  assign mac_24_5_reset = reset;
  assign mac_24_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_5_io_mulInput = mac_23_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_5_io_addInput = mac_24_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_6_clock = clock;
  assign mac_24_6_reset = reset;
  assign mac_24_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_6_io_mulInput = mac_23_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_6_io_addInput = mac_24_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_7_clock = clock;
  assign mac_24_7_reset = reset;
  assign mac_24_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_7_io_mulInput = mac_23_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_7_io_addInput = mac_24_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_8_clock = clock;
  assign mac_24_8_reset = reset;
  assign mac_24_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_8_io_mulInput = mac_23_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_8_io_addInput = mac_24_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_9_clock = clock;
  assign mac_24_9_reset = reset;
  assign mac_24_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_9_io_mulInput = mac_23_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_9_io_addInput = mac_24_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_10_clock = clock;
  assign mac_24_10_reset = reset;
  assign mac_24_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_10_io_mulInput = mac_23_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_10_io_addInput = mac_24_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_11_clock = clock;
  assign mac_24_11_reset = reset;
  assign mac_24_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_11_io_mulInput = mac_23_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_11_io_addInput = mac_24_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_12_clock = clock;
  assign mac_24_12_reset = reset;
  assign mac_24_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_12_io_mulInput = mac_23_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_12_io_addInput = mac_24_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_13_clock = clock;
  assign mac_24_13_reset = reset;
  assign mac_24_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_13_io_mulInput = mac_23_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_13_io_addInput = mac_24_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_14_clock = clock;
  assign mac_24_14_reset = reset;
  assign mac_24_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_14_io_mulInput = mac_23_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_14_io_addInput = mac_24_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_15_clock = clock;
  assign mac_24_15_reset = reset;
  assign mac_24_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_15_io_mulInput = mac_23_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_15_io_addInput = mac_24_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_16_clock = clock;
  assign mac_24_16_reset = reset;
  assign mac_24_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_16_io_mulInput = mac_23_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_16_io_addInput = mac_24_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_17_clock = clock;
  assign mac_24_17_reset = reset;
  assign mac_24_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_17_io_mulInput = mac_23_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_17_io_addInput = mac_24_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_18_clock = clock;
  assign mac_24_18_reset = reset;
  assign mac_24_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_18_io_mulInput = mac_23_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_18_io_addInput = mac_24_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_19_clock = clock;
  assign mac_24_19_reset = reset;
  assign mac_24_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_19_io_mulInput = mac_23_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_19_io_addInput = mac_24_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_20_clock = clock;
  assign mac_24_20_reset = reset;
  assign mac_24_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_20_io_mulInput = mac_23_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_20_io_addInput = mac_24_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_21_clock = clock;
  assign mac_24_21_reset = reset;
  assign mac_24_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_21_io_mulInput = mac_23_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_21_io_addInput = mac_24_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_22_clock = clock;
  assign mac_24_22_reset = reset;
  assign mac_24_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_22_io_mulInput = mac_23_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_22_io_addInput = mac_24_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_23_clock = clock;
  assign mac_24_23_reset = reset;
  assign mac_24_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_23_io_mulInput = mac_23_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_23_io_addInput = mac_24_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_24_clock = clock;
  assign mac_24_24_reset = reset;
  assign mac_24_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_24_io_mulInput = mac_23_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_24_io_addInput = mac_24_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_25_clock = clock;
  assign mac_24_25_reset = reset;
  assign mac_24_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_25_io_mulInput = mac_23_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_25_io_addInput = mac_24_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_26_clock = clock;
  assign mac_24_26_reset = reset;
  assign mac_24_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_26_io_mulInput = mac_23_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_26_io_addInput = mac_24_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_27_clock = clock;
  assign mac_24_27_reset = reset;
  assign mac_24_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_27_io_mulInput = mac_23_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_27_io_addInput = mac_24_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_28_clock = clock;
  assign mac_24_28_reset = reset;
  assign mac_24_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_28_io_mulInput = mac_23_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_28_io_addInput = mac_24_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_29_clock = clock;
  assign mac_24_29_reset = reset;
  assign mac_24_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_29_io_mulInput = mac_23_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_29_io_addInput = mac_24_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_30_clock = clock;
  assign mac_24_30_reset = reset;
  assign mac_24_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_30_io_mulInput = mac_23_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_30_io_addInput = mac_24_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_24_31_clock = clock;
  assign mac_24_31_reset = reset;
  assign mac_24_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_24_31_io_mulInput = mac_23_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_24_31_io_addInput = mac_24_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_0_clock = clock;
  assign mac_25_0_reset = reset;
  assign mac_25_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_25_0_io_mulInput = mac_24_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_25_0_io_addInput = bias_25; // @[InnerSystolicArray.scala 57:27]
  assign mac_25_1_clock = clock;
  assign mac_25_1_reset = reset;
  assign mac_25_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_1_io_mulInput = mac_24_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_1_io_addInput = mac_25_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_2_clock = clock;
  assign mac_25_2_reset = reset;
  assign mac_25_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_2_io_mulInput = mac_24_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_2_io_addInput = mac_25_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_3_clock = clock;
  assign mac_25_3_reset = reset;
  assign mac_25_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_3_io_mulInput = mac_24_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_3_io_addInput = mac_25_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_4_clock = clock;
  assign mac_25_4_reset = reset;
  assign mac_25_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_4_io_mulInput = mac_24_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_4_io_addInput = mac_25_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_5_clock = clock;
  assign mac_25_5_reset = reset;
  assign mac_25_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_5_io_mulInput = mac_24_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_5_io_addInput = mac_25_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_6_clock = clock;
  assign mac_25_6_reset = reset;
  assign mac_25_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_6_io_mulInput = mac_24_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_6_io_addInput = mac_25_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_7_clock = clock;
  assign mac_25_7_reset = reset;
  assign mac_25_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_7_io_mulInput = mac_24_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_7_io_addInput = mac_25_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_8_clock = clock;
  assign mac_25_8_reset = reset;
  assign mac_25_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_8_io_mulInput = mac_24_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_8_io_addInput = mac_25_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_9_clock = clock;
  assign mac_25_9_reset = reset;
  assign mac_25_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_9_io_mulInput = mac_24_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_9_io_addInput = mac_25_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_10_clock = clock;
  assign mac_25_10_reset = reset;
  assign mac_25_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_10_io_mulInput = mac_24_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_10_io_addInput = mac_25_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_11_clock = clock;
  assign mac_25_11_reset = reset;
  assign mac_25_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_11_io_mulInput = mac_24_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_11_io_addInput = mac_25_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_12_clock = clock;
  assign mac_25_12_reset = reset;
  assign mac_25_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_12_io_mulInput = mac_24_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_12_io_addInput = mac_25_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_13_clock = clock;
  assign mac_25_13_reset = reset;
  assign mac_25_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_13_io_mulInput = mac_24_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_13_io_addInput = mac_25_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_14_clock = clock;
  assign mac_25_14_reset = reset;
  assign mac_25_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_14_io_mulInput = mac_24_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_14_io_addInput = mac_25_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_15_clock = clock;
  assign mac_25_15_reset = reset;
  assign mac_25_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_15_io_mulInput = mac_24_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_15_io_addInput = mac_25_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_16_clock = clock;
  assign mac_25_16_reset = reset;
  assign mac_25_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_16_io_mulInput = mac_24_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_16_io_addInput = mac_25_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_17_clock = clock;
  assign mac_25_17_reset = reset;
  assign mac_25_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_17_io_mulInput = mac_24_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_17_io_addInput = mac_25_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_18_clock = clock;
  assign mac_25_18_reset = reset;
  assign mac_25_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_18_io_mulInput = mac_24_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_18_io_addInput = mac_25_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_19_clock = clock;
  assign mac_25_19_reset = reset;
  assign mac_25_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_19_io_mulInput = mac_24_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_19_io_addInput = mac_25_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_20_clock = clock;
  assign mac_25_20_reset = reset;
  assign mac_25_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_20_io_mulInput = mac_24_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_20_io_addInput = mac_25_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_21_clock = clock;
  assign mac_25_21_reset = reset;
  assign mac_25_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_21_io_mulInput = mac_24_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_21_io_addInput = mac_25_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_22_clock = clock;
  assign mac_25_22_reset = reset;
  assign mac_25_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_22_io_mulInput = mac_24_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_22_io_addInput = mac_25_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_23_clock = clock;
  assign mac_25_23_reset = reset;
  assign mac_25_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_23_io_mulInput = mac_24_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_23_io_addInput = mac_25_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_24_clock = clock;
  assign mac_25_24_reset = reset;
  assign mac_25_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_24_io_mulInput = mac_24_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_24_io_addInput = mac_25_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_25_clock = clock;
  assign mac_25_25_reset = reset;
  assign mac_25_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_25_io_mulInput = mac_24_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_25_io_addInput = mac_25_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_26_clock = clock;
  assign mac_25_26_reset = reset;
  assign mac_25_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_26_io_mulInput = mac_24_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_26_io_addInput = mac_25_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_27_clock = clock;
  assign mac_25_27_reset = reset;
  assign mac_25_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_27_io_mulInput = mac_24_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_27_io_addInput = mac_25_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_28_clock = clock;
  assign mac_25_28_reset = reset;
  assign mac_25_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_28_io_mulInput = mac_24_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_28_io_addInput = mac_25_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_29_clock = clock;
  assign mac_25_29_reset = reset;
  assign mac_25_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_29_io_mulInput = mac_24_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_29_io_addInput = mac_25_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_30_clock = clock;
  assign mac_25_30_reset = reset;
  assign mac_25_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_30_io_mulInput = mac_24_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_30_io_addInput = mac_25_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_25_31_clock = clock;
  assign mac_25_31_reset = reset;
  assign mac_25_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_25_31_io_mulInput = mac_24_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_25_31_io_addInput = mac_25_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_0_clock = clock;
  assign mac_26_0_reset = reset;
  assign mac_26_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_26_0_io_mulInput = mac_25_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_26_0_io_addInput = bias_26; // @[InnerSystolicArray.scala 57:27]
  assign mac_26_1_clock = clock;
  assign mac_26_1_reset = reset;
  assign mac_26_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_1_io_mulInput = mac_25_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_1_io_addInput = mac_26_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_2_clock = clock;
  assign mac_26_2_reset = reset;
  assign mac_26_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_2_io_mulInput = mac_25_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_2_io_addInput = mac_26_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_3_clock = clock;
  assign mac_26_3_reset = reset;
  assign mac_26_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_3_io_mulInput = mac_25_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_3_io_addInput = mac_26_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_4_clock = clock;
  assign mac_26_4_reset = reset;
  assign mac_26_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_4_io_mulInput = mac_25_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_4_io_addInput = mac_26_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_5_clock = clock;
  assign mac_26_5_reset = reset;
  assign mac_26_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_5_io_mulInput = mac_25_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_5_io_addInput = mac_26_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_6_clock = clock;
  assign mac_26_6_reset = reset;
  assign mac_26_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_6_io_mulInput = mac_25_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_6_io_addInput = mac_26_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_7_clock = clock;
  assign mac_26_7_reset = reset;
  assign mac_26_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_7_io_mulInput = mac_25_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_7_io_addInput = mac_26_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_8_clock = clock;
  assign mac_26_8_reset = reset;
  assign mac_26_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_8_io_mulInput = mac_25_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_8_io_addInput = mac_26_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_9_clock = clock;
  assign mac_26_9_reset = reset;
  assign mac_26_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_9_io_mulInput = mac_25_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_9_io_addInput = mac_26_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_10_clock = clock;
  assign mac_26_10_reset = reset;
  assign mac_26_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_10_io_mulInput = mac_25_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_10_io_addInput = mac_26_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_11_clock = clock;
  assign mac_26_11_reset = reset;
  assign mac_26_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_11_io_mulInput = mac_25_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_11_io_addInput = mac_26_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_12_clock = clock;
  assign mac_26_12_reset = reset;
  assign mac_26_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_12_io_mulInput = mac_25_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_12_io_addInput = mac_26_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_13_clock = clock;
  assign mac_26_13_reset = reset;
  assign mac_26_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_13_io_mulInput = mac_25_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_13_io_addInput = mac_26_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_14_clock = clock;
  assign mac_26_14_reset = reset;
  assign mac_26_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_14_io_mulInput = mac_25_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_14_io_addInput = mac_26_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_15_clock = clock;
  assign mac_26_15_reset = reset;
  assign mac_26_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_15_io_mulInput = mac_25_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_15_io_addInput = mac_26_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_16_clock = clock;
  assign mac_26_16_reset = reset;
  assign mac_26_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_16_io_mulInput = mac_25_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_16_io_addInput = mac_26_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_17_clock = clock;
  assign mac_26_17_reset = reset;
  assign mac_26_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_17_io_mulInput = mac_25_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_17_io_addInput = mac_26_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_18_clock = clock;
  assign mac_26_18_reset = reset;
  assign mac_26_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_18_io_mulInput = mac_25_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_18_io_addInput = mac_26_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_19_clock = clock;
  assign mac_26_19_reset = reset;
  assign mac_26_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_19_io_mulInput = mac_25_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_19_io_addInput = mac_26_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_20_clock = clock;
  assign mac_26_20_reset = reset;
  assign mac_26_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_20_io_mulInput = mac_25_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_20_io_addInput = mac_26_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_21_clock = clock;
  assign mac_26_21_reset = reset;
  assign mac_26_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_21_io_mulInput = mac_25_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_21_io_addInput = mac_26_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_22_clock = clock;
  assign mac_26_22_reset = reset;
  assign mac_26_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_22_io_mulInput = mac_25_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_22_io_addInput = mac_26_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_23_clock = clock;
  assign mac_26_23_reset = reset;
  assign mac_26_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_23_io_mulInput = mac_25_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_23_io_addInput = mac_26_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_24_clock = clock;
  assign mac_26_24_reset = reset;
  assign mac_26_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_24_io_mulInput = mac_25_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_24_io_addInput = mac_26_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_25_clock = clock;
  assign mac_26_25_reset = reset;
  assign mac_26_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_25_io_mulInput = mac_25_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_25_io_addInput = mac_26_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_26_clock = clock;
  assign mac_26_26_reset = reset;
  assign mac_26_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_26_io_mulInput = mac_25_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_26_io_addInput = mac_26_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_27_clock = clock;
  assign mac_26_27_reset = reset;
  assign mac_26_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_27_io_mulInput = mac_25_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_27_io_addInput = mac_26_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_28_clock = clock;
  assign mac_26_28_reset = reset;
  assign mac_26_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_28_io_mulInput = mac_25_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_28_io_addInput = mac_26_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_29_clock = clock;
  assign mac_26_29_reset = reset;
  assign mac_26_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_29_io_mulInput = mac_25_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_29_io_addInput = mac_26_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_30_clock = clock;
  assign mac_26_30_reset = reset;
  assign mac_26_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_30_io_mulInput = mac_25_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_30_io_addInput = mac_26_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_26_31_clock = clock;
  assign mac_26_31_reset = reset;
  assign mac_26_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_26_31_io_mulInput = mac_25_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_26_31_io_addInput = mac_26_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_0_clock = clock;
  assign mac_27_0_reset = reset;
  assign mac_27_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_27_0_io_mulInput = mac_26_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_27_0_io_addInput = bias_27; // @[InnerSystolicArray.scala 57:27]
  assign mac_27_1_clock = clock;
  assign mac_27_1_reset = reset;
  assign mac_27_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_1_io_mulInput = mac_26_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_1_io_addInput = mac_27_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_2_clock = clock;
  assign mac_27_2_reset = reset;
  assign mac_27_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_2_io_mulInput = mac_26_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_2_io_addInput = mac_27_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_3_clock = clock;
  assign mac_27_3_reset = reset;
  assign mac_27_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_3_io_mulInput = mac_26_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_3_io_addInput = mac_27_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_4_clock = clock;
  assign mac_27_4_reset = reset;
  assign mac_27_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_4_io_mulInput = mac_26_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_4_io_addInput = mac_27_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_5_clock = clock;
  assign mac_27_5_reset = reset;
  assign mac_27_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_5_io_mulInput = mac_26_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_5_io_addInput = mac_27_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_6_clock = clock;
  assign mac_27_6_reset = reset;
  assign mac_27_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_6_io_mulInput = mac_26_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_6_io_addInput = mac_27_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_7_clock = clock;
  assign mac_27_7_reset = reset;
  assign mac_27_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_7_io_mulInput = mac_26_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_7_io_addInput = mac_27_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_8_clock = clock;
  assign mac_27_8_reset = reset;
  assign mac_27_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_8_io_mulInput = mac_26_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_8_io_addInput = mac_27_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_9_clock = clock;
  assign mac_27_9_reset = reset;
  assign mac_27_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_9_io_mulInput = mac_26_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_9_io_addInput = mac_27_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_10_clock = clock;
  assign mac_27_10_reset = reset;
  assign mac_27_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_10_io_mulInput = mac_26_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_10_io_addInput = mac_27_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_11_clock = clock;
  assign mac_27_11_reset = reset;
  assign mac_27_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_11_io_mulInput = mac_26_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_11_io_addInput = mac_27_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_12_clock = clock;
  assign mac_27_12_reset = reset;
  assign mac_27_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_12_io_mulInput = mac_26_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_12_io_addInput = mac_27_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_13_clock = clock;
  assign mac_27_13_reset = reset;
  assign mac_27_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_13_io_mulInput = mac_26_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_13_io_addInput = mac_27_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_14_clock = clock;
  assign mac_27_14_reset = reset;
  assign mac_27_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_14_io_mulInput = mac_26_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_14_io_addInput = mac_27_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_15_clock = clock;
  assign mac_27_15_reset = reset;
  assign mac_27_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_15_io_mulInput = mac_26_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_15_io_addInput = mac_27_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_16_clock = clock;
  assign mac_27_16_reset = reset;
  assign mac_27_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_16_io_mulInput = mac_26_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_16_io_addInput = mac_27_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_17_clock = clock;
  assign mac_27_17_reset = reset;
  assign mac_27_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_17_io_mulInput = mac_26_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_17_io_addInput = mac_27_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_18_clock = clock;
  assign mac_27_18_reset = reset;
  assign mac_27_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_18_io_mulInput = mac_26_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_18_io_addInput = mac_27_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_19_clock = clock;
  assign mac_27_19_reset = reset;
  assign mac_27_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_19_io_mulInput = mac_26_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_19_io_addInput = mac_27_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_20_clock = clock;
  assign mac_27_20_reset = reset;
  assign mac_27_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_20_io_mulInput = mac_26_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_20_io_addInput = mac_27_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_21_clock = clock;
  assign mac_27_21_reset = reset;
  assign mac_27_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_21_io_mulInput = mac_26_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_21_io_addInput = mac_27_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_22_clock = clock;
  assign mac_27_22_reset = reset;
  assign mac_27_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_22_io_mulInput = mac_26_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_22_io_addInput = mac_27_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_23_clock = clock;
  assign mac_27_23_reset = reset;
  assign mac_27_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_23_io_mulInput = mac_26_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_23_io_addInput = mac_27_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_24_clock = clock;
  assign mac_27_24_reset = reset;
  assign mac_27_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_24_io_mulInput = mac_26_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_24_io_addInput = mac_27_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_25_clock = clock;
  assign mac_27_25_reset = reset;
  assign mac_27_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_25_io_mulInput = mac_26_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_25_io_addInput = mac_27_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_26_clock = clock;
  assign mac_27_26_reset = reset;
  assign mac_27_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_26_io_mulInput = mac_26_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_26_io_addInput = mac_27_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_27_clock = clock;
  assign mac_27_27_reset = reset;
  assign mac_27_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_27_io_mulInput = mac_26_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_27_io_addInput = mac_27_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_28_clock = clock;
  assign mac_27_28_reset = reset;
  assign mac_27_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_28_io_mulInput = mac_26_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_28_io_addInput = mac_27_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_29_clock = clock;
  assign mac_27_29_reset = reset;
  assign mac_27_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_29_io_mulInput = mac_26_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_29_io_addInput = mac_27_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_30_clock = clock;
  assign mac_27_30_reset = reset;
  assign mac_27_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_30_io_mulInput = mac_26_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_30_io_addInput = mac_27_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_27_31_clock = clock;
  assign mac_27_31_reset = reset;
  assign mac_27_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_27_31_io_mulInput = mac_26_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_27_31_io_addInput = mac_27_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_0_clock = clock;
  assign mac_28_0_reset = reset;
  assign mac_28_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_28_0_io_mulInput = mac_27_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_28_0_io_addInput = bias_28; // @[InnerSystolicArray.scala 57:27]
  assign mac_28_1_clock = clock;
  assign mac_28_1_reset = reset;
  assign mac_28_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_1_io_mulInput = mac_27_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_1_io_addInput = mac_28_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_2_clock = clock;
  assign mac_28_2_reset = reset;
  assign mac_28_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_2_io_mulInput = mac_27_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_2_io_addInput = mac_28_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_3_clock = clock;
  assign mac_28_3_reset = reset;
  assign mac_28_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_3_io_mulInput = mac_27_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_3_io_addInput = mac_28_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_4_clock = clock;
  assign mac_28_4_reset = reset;
  assign mac_28_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_4_io_mulInput = mac_27_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_4_io_addInput = mac_28_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_5_clock = clock;
  assign mac_28_5_reset = reset;
  assign mac_28_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_5_io_mulInput = mac_27_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_5_io_addInput = mac_28_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_6_clock = clock;
  assign mac_28_6_reset = reset;
  assign mac_28_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_6_io_mulInput = mac_27_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_6_io_addInput = mac_28_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_7_clock = clock;
  assign mac_28_7_reset = reset;
  assign mac_28_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_7_io_mulInput = mac_27_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_7_io_addInput = mac_28_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_8_clock = clock;
  assign mac_28_8_reset = reset;
  assign mac_28_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_8_io_mulInput = mac_27_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_8_io_addInput = mac_28_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_9_clock = clock;
  assign mac_28_9_reset = reset;
  assign mac_28_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_9_io_mulInput = mac_27_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_9_io_addInput = mac_28_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_10_clock = clock;
  assign mac_28_10_reset = reset;
  assign mac_28_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_10_io_mulInput = mac_27_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_10_io_addInput = mac_28_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_11_clock = clock;
  assign mac_28_11_reset = reset;
  assign mac_28_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_11_io_mulInput = mac_27_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_11_io_addInput = mac_28_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_12_clock = clock;
  assign mac_28_12_reset = reset;
  assign mac_28_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_12_io_mulInput = mac_27_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_12_io_addInput = mac_28_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_13_clock = clock;
  assign mac_28_13_reset = reset;
  assign mac_28_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_13_io_mulInput = mac_27_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_13_io_addInput = mac_28_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_14_clock = clock;
  assign mac_28_14_reset = reset;
  assign mac_28_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_14_io_mulInput = mac_27_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_14_io_addInput = mac_28_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_15_clock = clock;
  assign mac_28_15_reset = reset;
  assign mac_28_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_15_io_mulInput = mac_27_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_15_io_addInput = mac_28_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_16_clock = clock;
  assign mac_28_16_reset = reset;
  assign mac_28_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_16_io_mulInput = mac_27_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_16_io_addInput = mac_28_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_17_clock = clock;
  assign mac_28_17_reset = reset;
  assign mac_28_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_17_io_mulInput = mac_27_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_17_io_addInput = mac_28_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_18_clock = clock;
  assign mac_28_18_reset = reset;
  assign mac_28_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_18_io_mulInput = mac_27_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_18_io_addInput = mac_28_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_19_clock = clock;
  assign mac_28_19_reset = reset;
  assign mac_28_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_19_io_mulInput = mac_27_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_19_io_addInput = mac_28_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_20_clock = clock;
  assign mac_28_20_reset = reset;
  assign mac_28_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_20_io_mulInput = mac_27_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_20_io_addInput = mac_28_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_21_clock = clock;
  assign mac_28_21_reset = reset;
  assign mac_28_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_21_io_mulInput = mac_27_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_21_io_addInput = mac_28_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_22_clock = clock;
  assign mac_28_22_reset = reset;
  assign mac_28_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_22_io_mulInput = mac_27_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_22_io_addInput = mac_28_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_23_clock = clock;
  assign mac_28_23_reset = reset;
  assign mac_28_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_23_io_mulInput = mac_27_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_23_io_addInput = mac_28_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_24_clock = clock;
  assign mac_28_24_reset = reset;
  assign mac_28_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_24_io_mulInput = mac_27_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_24_io_addInput = mac_28_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_25_clock = clock;
  assign mac_28_25_reset = reset;
  assign mac_28_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_25_io_mulInput = mac_27_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_25_io_addInput = mac_28_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_26_clock = clock;
  assign mac_28_26_reset = reset;
  assign mac_28_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_26_io_mulInput = mac_27_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_26_io_addInput = mac_28_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_27_clock = clock;
  assign mac_28_27_reset = reset;
  assign mac_28_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_27_io_mulInput = mac_27_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_27_io_addInput = mac_28_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_28_clock = clock;
  assign mac_28_28_reset = reset;
  assign mac_28_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_28_io_mulInput = mac_27_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_28_io_addInput = mac_28_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_29_clock = clock;
  assign mac_28_29_reset = reset;
  assign mac_28_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_29_io_mulInput = mac_27_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_29_io_addInput = mac_28_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_30_clock = clock;
  assign mac_28_30_reset = reset;
  assign mac_28_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_30_io_mulInput = mac_27_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_30_io_addInput = mac_28_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_28_31_clock = clock;
  assign mac_28_31_reset = reset;
  assign mac_28_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_28_31_io_mulInput = mac_27_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_28_31_io_addInput = mac_28_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_0_clock = clock;
  assign mac_29_0_reset = reset;
  assign mac_29_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_29_0_io_mulInput = mac_28_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_29_0_io_addInput = bias_29; // @[InnerSystolicArray.scala 57:27]
  assign mac_29_1_clock = clock;
  assign mac_29_1_reset = reset;
  assign mac_29_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_1_io_mulInput = mac_28_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_1_io_addInput = mac_29_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_2_clock = clock;
  assign mac_29_2_reset = reset;
  assign mac_29_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_2_io_mulInput = mac_28_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_2_io_addInput = mac_29_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_3_clock = clock;
  assign mac_29_3_reset = reset;
  assign mac_29_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_3_io_mulInput = mac_28_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_3_io_addInput = mac_29_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_4_clock = clock;
  assign mac_29_4_reset = reset;
  assign mac_29_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_4_io_mulInput = mac_28_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_4_io_addInput = mac_29_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_5_clock = clock;
  assign mac_29_5_reset = reset;
  assign mac_29_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_5_io_mulInput = mac_28_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_5_io_addInput = mac_29_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_6_clock = clock;
  assign mac_29_6_reset = reset;
  assign mac_29_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_6_io_mulInput = mac_28_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_6_io_addInput = mac_29_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_7_clock = clock;
  assign mac_29_7_reset = reset;
  assign mac_29_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_7_io_mulInput = mac_28_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_7_io_addInput = mac_29_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_8_clock = clock;
  assign mac_29_8_reset = reset;
  assign mac_29_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_8_io_mulInput = mac_28_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_8_io_addInput = mac_29_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_9_clock = clock;
  assign mac_29_9_reset = reset;
  assign mac_29_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_9_io_mulInput = mac_28_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_9_io_addInput = mac_29_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_10_clock = clock;
  assign mac_29_10_reset = reset;
  assign mac_29_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_10_io_mulInput = mac_28_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_10_io_addInput = mac_29_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_11_clock = clock;
  assign mac_29_11_reset = reset;
  assign mac_29_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_11_io_mulInput = mac_28_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_11_io_addInput = mac_29_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_12_clock = clock;
  assign mac_29_12_reset = reset;
  assign mac_29_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_12_io_mulInput = mac_28_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_12_io_addInput = mac_29_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_13_clock = clock;
  assign mac_29_13_reset = reset;
  assign mac_29_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_13_io_mulInput = mac_28_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_13_io_addInput = mac_29_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_14_clock = clock;
  assign mac_29_14_reset = reset;
  assign mac_29_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_14_io_mulInput = mac_28_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_14_io_addInput = mac_29_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_15_clock = clock;
  assign mac_29_15_reset = reset;
  assign mac_29_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_15_io_mulInput = mac_28_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_15_io_addInput = mac_29_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_16_clock = clock;
  assign mac_29_16_reset = reset;
  assign mac_29_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_16_io_mulInput = mac_28_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_16_io_addInput = mac_29_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_17_clock = clock;
  assign mac_29_17_reset = reset;
  assign mac_29_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_17_io_mulInput = mac_28_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_17_io_addInput = mac_29_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_18_clock = clock;
  assign mac_29_18_reset = reset;
  assign mac_29_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_18_io_mulInput = mac_28_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_18_io_addInput = mac_29_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_19_clock = clock;
  assign mac_29_19_reset = reset;
  assign mac_29_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_19_io_mulInput = mac_28_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_19_io_addInput = mac_29_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_20_clock = clock;
  assign mac_29_20_reset = reset;
  assign mac_29_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_20_io_mulInput = mac_28_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_20_io_addInput = mac_29_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_21_clock = clock;
  assign mac_29_21_reset = reset;
  assign mac_29_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_21_io_mulInput = mac_28_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_21_io_addInput = mac_29_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_22_clock = clock;
  assign mac_29_22_reset = reset;
  assign mac_29_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_22_io_mulInput = mac_28_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_22_io_addInput = mac_29_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_23_clock = clock;
  assign mac_29_23_reset = reset;
  assign mac_29_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_23_io_mulInput = mac_28_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_23_io_addInput = mac_29_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_24_clock = clock;
  assign mac_29_24_reset = reset;
  assign mac_29_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_24_io_mulInput = mac_28_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_24_io_addInput = mac_29_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_25_clock = clock;
  assign mac_29_25_reset = reset;
  assign mac_29_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_25_io_mulInput = mac_28_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_25_io_addInput = mac_29_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_26_clock = clock;
  assign mac_29_26_reset = reset;
  assign mac_29_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_26_io_mulInput = mac_28_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_26_io_addInput = mac_29_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_27_clock = clock;
  assign mac_29_27_reset = reset;
  assign mac_29_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_27_io_mulInput = mac_28_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_27_io_addInput = mac_29_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_28_clock = clock;
  assign mac_29_28_reset = reset;
  assign mac_29_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_28_io_mulInput = mac_28_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_28_io_addInput = mac_29_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_29_clock = clock;
  assign mac_29_29_reset = reset;
  assign mac_29_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_29_io_mulInput = mac_28_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_29_io_addInput = mac_29_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_30_clock = clock;
  assign mac_29_30_reset = reset;
  assign mac_29_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_30_io_mulInput = mac_28_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_30_io_addInput = mac_29_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_29_31_clock = clock;
  assign mac_29_31_reset = reset;
  assign mac_29_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_29_31_io_mulInput = mac_28_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_29_31_io_addInput = mac_29_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_0_clock = clock;
  assign mac_30_0_reset = reset;
  assign mac_30_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_30_0_io_mulInput = mac_29_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_30_0_io_addInput = bias_30; // @[InnerSystolicArray.scala 57:27]
  assign mac_30_1_clock = clock;
  assign mac_30_1_reset = reset;
  assign mac_30_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_1_io_mulInput = mac_29_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_1_io_addInput = mac_30_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_2_clock = clock;
  assign mac_30_2_reset = reset;
  assign mac_30_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_2_io_mulInput = mac_29_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_2_io_addInput = mac_30_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_3_clock = clock;
  assign mac_30_3_reset = reset;
  assign mac_30_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_3_io_mulInput = mac_29_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_3_io_addInput = mac_30_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_4_clock = clock;
  assign mac_30_4_reset = reset;
  assign mac_30_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_4_io_mulInput = mac_29_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_4_io_addInput = mac_30_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_5_clock = clock;
  assign mac_30_5_reset = reset;
  assign mac_30_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_5_io_mulInput = mac_29_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_5_io_addInput = mac_30_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_6_clock = clock;
  assign mac_30_6_reset = reset;
  assign mac_30_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_6_io_mulInput = mac_29_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_6_io_addInput = mac_30_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_7_clock = clock;
  assign mac_30_7_reset = reset;
  assign mac_30_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_7_io_mulInput = mac_29_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_7_io_addInput = mac_30_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_8_clock = clock;
  assign mac_30_8_reset = reset;
  assign mac_30_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_8_io_mulInput = mac_29_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_8_io_addInput = mac_30_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_9_clock = clock;
  assign mac_30_9_reset = reset;
  assign mac_30_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_9_io_mulInput = mac_29_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_9_io_addInput = mac_30_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_10_clock = clock;
  assign mac_30_10_reset = reset;
  assign mac_30_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_10_io_mulInput = mac_29_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_10_io_addInput = mac_30_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_11_clock = clock;
  assign mac_30_11_reset = reset;
  assign mac_30_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_11_io_mulInput = mac_29_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_11_io_addInput = mac_30_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_12_clock = clock;
  assign mac_30_12_reset = reset;
  assign mac_30_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_12_io_mulInput = mac_29_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_12_io_addInput = mac_30_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_13_clock = clock;
  assign mac_30_13_reset = reset;
  assign mac_30_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_13_io_mulInput = mac_29_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_13_io_addInput = mac_30_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_14_clock = clock;
  assign mac_30_14_reset = reset;
  assign mac_30_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_14_io_mulInput = mac_29_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_14_io_addInput = mac_30_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_15_clock = clock;
  assign mac_30_15_reset = reset;
  assign mac_30_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_15_io_mulInput = mac_29_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_15_io_addInput = mac_30_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_16_clock = clock;
  assign mac_30_16_reset = reset;
  assign mac_30_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_16_io_mulInput = mac_29_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_16_io_addInput = mac_30_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_17_clock = clock;
  assign mac_30_17_reset = reset;
  assign mac_30_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_17_io_mulInput = mac_29_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_17_io_addInput = mac_30_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_18_clock = clock;
  assign mac_30_18_reset = reset;
  assign mac_30_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_18_io_mulInput = mac_29_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_18_io_addInput = mac_30_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_19_clock = clock;
  assign mac_30_19_reset = reset;
  assign mac_30_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_19_io_mulInput = mac_29_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_19_io_addInput = mac_30_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_20_clock = clock;
  assign mac_30_20_reset = reset;
  assign mac_30_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_20_io_mulInput = mac_29_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_20_io_addInput = mac_30_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_21_clock = clock;
  assign mac_30_21_reset = reset;
  assign mac_30_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_21_io_mulInput = mac_29_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_21_io_addInput = mac_30_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_22_clock = clock;
  assign mac_30_22_reset = reset;
  assign mac_30_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_22_io_mulInput = mac_29_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_22_io_addInput = mac_30_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_23_clock = clock;
  assign mac_30_23_reset = reset;
  assign mac_30_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_23_io_mulInput = mac_29_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_23_io_addInput = mac_30_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_24_clock = clock;
  assign mac_30_24_reset = reset;
  assign mac_30_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_24_io_mulInput = mac_29_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_24_io_addInput = mac_30_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_25_clock = clock;
  assign mac_30_25_reset = reset;
  assign mac_30_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_25_io_mulInput = mac_29_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_25_io_addInput = mac_30_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_26_clock = clock;
  assign mac_30_26_reset = reset;
  assign mac_30_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_26_io_mulInput = mac_29_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_26_io_addInput = mac_30_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_27_clock = clock;
  assign mac_30_27_reset = reset;
  assign mac_30_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_27_io_mulInput = mac_29_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_27_io_addInput = mac_30_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_28_clock = clock;
  assign mac_30_28_reset = reset;
  assign mac_30_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_28_io_mulInput = mac_29_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_28_io_addInput = mac_30_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_29_clock = clock;
  assign mac_30_29_reset = reset;
  assign mac_30_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_29_io_mulInput = mac_29_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_29_io_addInput = mac_30_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_30_clock = clock;
  assign mac_30_30_reset = reset;
  assign mac_30_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_30_io_mulInput = mac_29_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_30_io_addInput = mac_30_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_30_31_clock = clock;
  assign mac_30_31_reset = reset;
  assign mac_30_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_30_31_io_mulInput = mac_29_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_30_31_io_addInput = mac_30_30_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_0_clock = clock;
  assign mac_31_0_reset = reset;
  assign mac_31_0_io_load = io_load; // @[InnerSystolicArray.scala 60:25]
  assign mac_31_0_io_mulInput = mac_30_0_io_passthrough; // @[InnerSystolicArray.scala 59:29]
  assign mac_31_0_io_addInput = bias_31; // @[InnerSystolicArray.scala 57:27]
  assign mac_31_1_clock = clock;
  assign mac_31_1_reset = reset;
  assign mac_31_1_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_1_io_mulInput = mac_30_1_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_1_io_addInput = mac_31_0_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_2_clock = clock;
  assign mac_31_2_reset = reset;
  assign mac_31_2_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_2_io_mulInput = mac_30_2_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_2_io_addInput = mac_31_1_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_3_clock = clock;
  assign mac_31_3_reset = reset;
  assign mac_31_3_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_3_io_mulInput = mac_30_3_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_3_io_addInput = mac_31_2_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_4_clock = clock;
  assign mac_31_4_reset = reset;
  assign mac_31_4_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_4_io_mulInput = mac_30_4_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_4_io_addInput = mac_31_3_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_5_clock = clock;
  assign mac_31_5_reset = reset;
  assign mac_31_5_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_5_io_mulInput = mac_30_5_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_5_io_addInput = mac_31_4_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_6_clock = clock;
  assign mac_31_6_reset = reset;
  assign mac_31_6_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_6_io_mulInput = mac_30_6_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_6_io_addInput = mac_31_5_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_7_clock = clock;
  assign mac_31_7_reset = reset;
  assign mac_31_7_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_7_io_mulInput = mac_30_7_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_7_io_addInput = mac_31_6_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_8_clock = clock;
  assign mac_31_8_reset = reset;
  assign mac_31_8_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_8_io_mulInput = mac_30_8_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_8_io_addInput = mac_31_7_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_9_clock = clock;
  assign mac_31_9_reset = reset;
  assign mac_31_9_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_9_io_mulInput = mac_30_9_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_9_io_addInput = mac_31_8_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_10_clock = clock;
  assign mac_31_10_reset = reset;
  assign mac_31_10_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_10_io_mulInput = mac_30_10_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_10_io_addInput = mac_31_9_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_11_clock = clock;
  assign mac_31_11_reset = reset;
  assign mac_31_11_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_11_io_mulInput = mac_30_11_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_11_io_addInput = mac_31_10_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_12_clock = clock;
  assign mac_31_12_reset = reset;
  assign mac_31_12_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_12_io_mulInput = mac_30_12_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_12_io_addInput = mac_31_11_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_13_clock = clock;
  assign mac_31_13_reset = reset;
  assign mac_31_13_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_13_io_mulInput = mac_30_13_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_13_io_addInput = mac_31_12_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_14_clock = clock;
  assign mac_31_14_reset = reset;
  assign mac_31_14_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_14_io_mulInput = mac_30_14_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_14_io_addInput = mac_31_13_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_15_clock = clock;
  assign mac_31_15_reset = reset;
  assign mac_31_15_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_15_io_mulInput = mac_30_15_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_15_io_addInput = mac_31_14_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_16_clock = clock;
  assign mac_31_16_reset = reset;
  assign mac_31_16_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_16_io_mulInput = mac_30_16_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_16_io_addInput = mac_31_15_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_17_clock = clock;
  assign mac_31_17_reset = reset;
  assign mac_31_17_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_17_io_mulInput = mac_30_17_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_17_io_addInput = mac_31_16_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_18_clock = clock;
  assign mac_31_18_reset = reset;
  assign mac_31_18_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_18_io_mulInput = mac_30_18_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_18_io_addInput = mac_31_17_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_19_clock = clock;
  assign mac_31_19_reset = reset;
  assign mac_31_19_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_19_io_mulInput = mac_30_19_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_19_io_addInput = mac_31_18_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_20_clock = clock;
  assign mac_31_20_reset = reset;
  assign mac_31_20_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_20_io_mulInput = mac_30_20_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_20_io_addInput = mac_31_19_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_21_clock = clock;
  assign mac_31_21_reset = reset;
  assign mac_31_21_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_21_io_mulInput = mac_30_21_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_21_io_addInput = mac_31_20_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_22_clock = clock;
  assign mac_31_22_reset = reset;
  assign mac_31_22_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_22_io_mulInput = mac_30_22_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_22_io_addInput = mac_31_21_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_23_clock = clock;
  assign mac_31_23_reset = reset;
  assign mac_31_23_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_23_io_mulInput = mac_30_23_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_23_io_addInput = mac_31_22_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_24_clock = clock;
  assign mac_31_24_reset = reset;
  assign mac_31_24_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_24_io_mulInput = mac_30_24_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_24_io_addInput = mac_31_23_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_25_clock = clock;
  assign mac_31_25_reset = reset;
  assign mac_31_25_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_25_io_mulInput = mac_30_25_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_25_io_addInput = mac_31_24_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_26_clock = clock;
  assign mac_31_26_reset = reset;
  assign mac_31_26_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_26_io_mulInput = mac_30_26_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_26_io_addInput = mac_31_25_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_27_clock = clock;
  assign mac_31_27_reset = reset;
  assign mac_31_27_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_27_io_mulInput = mac_30_27_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_27_io_addInput = mac_31_26_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_28_clock = clock;
  assign mac_31_28_reset = reset;
  assign mac_31_28_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_28_io_mulInput = mac_30_28_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_28_io_addInput = mac_31_27_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_29_clock = clock;
  assign mac_31_29_reset = reset;
  assign mac_31_29_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_29_io_mulInput = mac_30_29_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_29_io_addInput = mac_31_28_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_30_clock = clock;
  assign mac_31_30_reset = reset;
  assign mac_31_30_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_30_io_mulInput = mac_30_30_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_30_io_addInput = mac_31_29_io_output; // @[InnerSystolicArray.scala 68:29]
  assign mac_31_31_clock = clock;
  assign mac_31_31_reset = reset;
  assign mac_31_31_io_load = io_load; // @[InnerSystolicArray.scala 69:25]
  assign mac_31_31_io_mulInput = mac_30_31_io_passthrough; // @[InnerSystolicArray.scala 67:29]
  assign mac_31_31_io_addInput = mac_31_30_io_output; // @[InnerSystolicArray.scala 68:29]
  always @(posedge clock) begin
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_0 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_0 <= io_weight_0; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_1 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_1 <= io_weight_1; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_2 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_2 <= io_weight_2; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_3 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_3 <= io_weight_3; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_4 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_4 <= io_weight_4; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_5 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_5 <= io_weight_5; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_6 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_6 <= io_weight_6; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_7 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_7 <= io_weight_7; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_8 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_8 <= io_weight_8; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_9 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_9 <= io_weight_9; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_10 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_10 <= io_weight_10; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_11 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_11 <= io_weight_11; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_12 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_12 <= io_weight_12; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_13 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_13 <= io_weight_13; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_14 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_14 <= io_weight_14; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_15 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_15 <= io_weight_15; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_16 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_16 <= io_weight_16; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_17 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_17 <= io_weight_17; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_18 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_18 <= io_weight_18; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_19 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_19 <= io_weight_19; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_20 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_20 <= io_weight_20; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_21 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_21 <= io_weight_21; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_22 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_22 <= io_weight_22; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_23 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_23 <= io_weight_23; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_24 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_24 <= io_weight_24; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_25 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_25 <= io_weight_25; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_26 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_26 <= io_weight_26; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_27 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_27 <= io_weight_27; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_28 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_28 <= io_weight_28; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_29 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_29 <= io_weight_29; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_30 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_30 <= io_weight_30; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[InnerSystolicArray.scala 37:20]
      bias_31 <= 16'sh0; // @[InnerSystolicArray.scala 37:20]
    end else if (io_load) begin // @[InnerSystolicArray.scala 38:19]
      bias_31 <= io_weight_31; // @[InnerSystolicArray.scala 39:9]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_1_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_1_io_mulInput_sr_0 <= io_input_1; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_2_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_2_io_mulInput_sr_0 <= io_input_2; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_2_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_2_io_mulInput_sr_1 <= mac_0_2_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_3_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_3_io_mulInput_sr_0 <= io_input_3; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_3_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_3_io_mulInput_sr_1 <= mac_0_3_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_3_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_3_io_mulInput_sr_2 <= mac_0_3_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_4_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_4_io_mulInput_sr_0 <= io_input_4; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_4_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_4_io_mulInput_sr_1 <= mac_0_4_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_4_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_4_io_mulInput_sr_2 <= mac_0_4_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_4_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_4_io_mulInput_sr_3 <= mac_0_4_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_5_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_5_io_mulInput_sr_0 <= io_input_5; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_5_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_5_io_mulInput_sr_1 <= mac_0_5_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_5_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_5_io_mulInput_sr_2 <= mac_0_5_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_5_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_5_io_mulInput_sr_3 <= mac_0_5_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_5_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_5_io_mulInput_sr_4 <= mac_0_5_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_6_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_6_io_mulInput_sr_0 <= io_input_6; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_6_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_6_io_mulInput_sr_1 <= mac_0_6_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_6_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_6_io_mulInput_sr_2 <= mac_0_6_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_6_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_6_io_mulInput_sr_3 <= mac_0_6_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_6_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_6_io_mulInput_sr_4 <= mac_0_6_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_6_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_6_io_mulInput_sr_5 <= mac_0_6_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_7_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_7_io_mulInput_sr_0 <= io_input_7; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_7_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_7_io_mulInput_sr_1 <= mac_0_7_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_7_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_7_io_mulInput_sr_2 <= mac_0_7_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_7_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_7_io_mulInput_sr_3 <= mac_0_7_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_7_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_7_io_mulInput_sr_4 <= mac_0_7_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_7_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_7_io_mulInput_sr_5 <= mac_0_7_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_7_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_7_io_mulInput_sr_6 <= mac_0_7_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_8_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_8_io_mulInput_sr_0 <= io_input_8; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_8_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_8_io_mulInput_sr_1 <= mac_0_8_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_8_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_8_io_mulInput_sr_2 <= mac_0_8_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_8_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_8_io_mulInput_sr_3 <= mac_0_8_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_8_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_8_io_mulInput_sr_4 <= mac_0_8_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_8_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_8_io_mulInput_sr_5 <= mac_0_8_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_8_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_8_io_mulInput_sr_6 <= mac_0_8_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_8_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_8_io_mulInput_sr_7 <= mac_0_8_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_9_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_9_io_mulInput_sr_0 <= io_input_9; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_9_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_9_io_mulInput_sr_1 <= mac_0_9_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_9_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_9_io_mulInput_sr_2 <= mac_0_9_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_9_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_9_io_mulInput_sr_3 <= mac_0_9_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_9_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_9_io_mulInput_sr_4 <= mac_0_9_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_9_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_9_io_mulInput_sr_5 <= mac_0_9_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_9_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_9_io_mulInput_sr_6 <= mac_0_9_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_9_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_9_io_mulInput_sr_7 <= mac_0_9_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_9_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_9_io_mulInput_sr_8 <= mac_0_9_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_10_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_10_io_mulInput_sr_0 <= io_input_10; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_10_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_10_io_mulInput_sr_1 <= mac_0_10_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_10_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_10_io_mulInput_sr_2 <= mac_0_10_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_10_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_10_io_mulInput_sr_3 <= mac_0_10_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_10_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_10_io_mulInput_sr_4 <= mac_0_10_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_10_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_10_io_mulInput_sr_5 <= mac_0_10_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_10_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_10_io_mulInput_sr_6 <= mac_0_10_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_10_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_10_io_mulInput_sr_7 <= mac_0_10_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_10_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_10_io_mulInput_sr_8 <= mac_0_10_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_10_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_10_io_mulInput_sr_9 <= mac_0_10_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_0 <= io_input_11; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_1 <= mac_0_11_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_2 <= mac_0_11_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_3 <= mac_0_11_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_4 <= mac_0_11_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_5 <= mac_0_11_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_6 <= mac_0_11_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_7 <= mac_0_11_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_8 <= mac_0_11_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_9 <= mac_0_11_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_11_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_11_io_mulInput_sr_10 <= mac_0_11_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_0 <= io_input_12; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_1 <= mac_0_12_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_2 <= mac_0_12_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_3 <= mac_0_12_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_4 <= mac_0_12_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_5 <= mac_0_12_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_6 <= mac_0_12_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_7 <= mac_0_12_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_8 <= mac_0_12_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_9 <= mac_0_12_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_10 <= mac_0_12_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_12_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_12_io_mulInput_sr_11 <= mac_0_12_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_0 <= io_input_13; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_1 <= mac_0_13_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_2 <= mac_0_13_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_3 <= mac_0_13_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_4 <= mac_0_13_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_5 <= mac_0_13_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_6 <= mac_0_13_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_7 <= mac_0_13_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_8 <= mac_0_13_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_9 <= mac_0_13_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_10 <= mac_0_13_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_11 <= mac_0_13_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_13_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_13_io_mulInput_sr_12 <= mac_0_13_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_0 <= io_input_14; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_1 <= mac_0_14_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_2 <= mac_0_14_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_3 <= mac_0_14_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_4 <= mac_0_14_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_5 <= mac_0_14_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_6 <= mac_0_14_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_7 <= mac_0_14_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_8 <= mac_0_14_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_9 <= mac_0_14_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_10 <= mac_0_14_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_11 <= mac_0_14_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_12 <= mac_0_14_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_14_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_14_io_mulInput_sr_13 <= mac_0_14_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_0 <= io_input_15; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_1 <= mac_0_15_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_2 <= mac_0_15_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_3 <= mac_0_15_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_4 <= mac_0_15_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_5 <= mac_0_15_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_6 <= mac_0_15_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_7 <= mac_0_15_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_8 <= mac_0_15_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_9 <= mac_0_15_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_10 <= mac_0_15_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_11 <= mac_0_15_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_12 <= mac_0_15_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_13 <= mac_0_15_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_15_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_15_io_mulInput_sr_14 <= mac_0_15_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_0 <= io_input_16; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_1 <= mac_0_16_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_2 <= mac_0_16_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_3 <= mac_0_16_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_4 <= mac_0_16_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_5 <= mac_0_16_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_6 <= mac_0_16_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_7 <= mac_0_16_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_8 <= mac_0_16_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_9 <= mac_0_16_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_10 <= mac_0_16_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_11 <= mac_0_16_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_12 <= mac_0_16_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_13 <= mac_0_16_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_14 <= mac_0_16_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_16_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_16_io_mulInput_sr_15 <= mac_0_16_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_0 <= io_input_17; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_1 <= mac_0_17_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_2 <= mac_0_17_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_3 <= mac_0_17_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_4 <= mac_0_17_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_5 <= mac_0_17_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_6 <= mac_0_17_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_7 <= mac_0_17_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_8 <= mac_0_17_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_9 <= mac_0_17_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_10 <= mac_0_17_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_11 <= mac_0_17_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_12 <= mac_0_17_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_13 <= mac_0_17_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_14 <= mac_0_17_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_15 <= mac_0_17_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_17_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_17_io_mulInput_sr_16 <= mac_0_17_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_0 <= io_input_18; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_1 <= mac_0_18_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_2 <= mac_0_18_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_3 <= mac_0_18_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_4 <= mac_0_18_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_5 <= mac_0_18_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_6 <= mac_0_18_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_7 <= mac_0_18_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_8 <= mac_0_18_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_9 <= mac_0_18_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_10 <= mac_0_18_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_11 <= mac_0_18_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_12 <= mac_0_18_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_13 <= mac_0_18_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_14 <= mac_0_18_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_15 <= mac_0_18_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_16 <= mac_0_18_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_18_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_18_io_mulInput_sr_17 <= mac_0_18_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_0 <= io_input_19; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_1 <= mac_0_19_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_2 <= mac_0_19_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_3 <= mac_0_19_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_4 <= mac_0_19_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_5 <= mac_0_19_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_6 <= mac_0_19_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_7 <= mac_0_19_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_8 <= mac_0_19_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_9 <= mac_0_19_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_10 <= mac_0_19_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_11 <= mac_0_19_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_12 <= mac_0_19_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_13 <= mac_0_19_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_14 <= mac_0_19_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_15 <= mac_0_19_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_16 <= mac_0_19_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_17 <= mac_0_19_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_19_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_19_io_mulInput_sr_18 <= mac_0_19_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_0 <= io_input_20; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_1 <= mac_0_20_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_2 <= mac_0_20_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_3 <= mac_0_20_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_4 <= mac_0_20_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_5 <= mac_0_20_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_6 <= mac_0_20_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_7 <= mac_0_20_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_8 <= mac_0_20_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_9 <= mac_0_20_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_10 <= mac_0_20_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_11 <= mac_0_20_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_12 <= mac_0_20_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_13 <= mac_0_20_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_14 <= mac_0_20_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_15 <= mac_0_20_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_16 <= mac_0_20_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_17 <= mac_0_20_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_18 <= mac_0_20_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_20_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_20_io_mulInput_sr_19 <= mac_0_20_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_0 <= io_input_21; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_1 <= mac_0_21_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_2 <= mac_0_21_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_3 <= mac_0_21_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_4 <= mac_0_21_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_5 <= mac_0_21_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_6 <= mac_0_21_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_7 <= mac_0_21_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_8 <= mac_0_21_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_9 <= mac_0_21_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_10 <= mac_0_21_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_11 <= mac_0_21_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_12 <= mac_0_21_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_13 <= mac_0_21_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_14 <= mac_0_21_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_15 <= mac_0_21_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_16 <= mac_0_21_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_17 <= mac_0_21_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_18 <= mac_0_21_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_19 <= mac_0_21_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_21_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_21_io_mulInput_sr_20 <= mac_0_21_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_0 <= io_input_22; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_1 <= mac_0_22_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_2 <= mac_0_22_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_3 <= mac_0_22_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_4 <= mac_0_22_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_5 <= mac_0_22_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_6 <= mac_0_22_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_7 <= mac_0_22_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_8 <= mac_0_22_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_9 <= mac_0_22_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_10 <= mac_0_22_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_11 <= mac_0_22_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_12 <= mac_0_22_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_13 <= mac_0_22_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_14 <= mac_0_22_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_15 <= mac_0_22_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_16 <= mac_0_22_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_17 <= mac_0_22_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_18 <= mac_0_22_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_19 <= mac_0_22_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_20 <= mac_0_22_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_22_io_mulInput_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_22_io_mulInput_sr_21 <= mac_0_22_io_mulInput_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_0 <= io_input_23; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_1 <= mac_0_23_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_2 <= mac_0_23_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_3 <= mac_0_23_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_4 <= mac_0_23_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_5 <= mac_0_23_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_6 <= mac_0_23_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_7 <= mac_0_23_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_8 <= mac_0_23_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_9 <= mac_0_23_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_10 <= mac_0_23_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_11 <= mac_0_23_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_12 <= mac_0_23_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_13 <= mac_0_23_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_14 <= mac_0_23_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_15 <= mac_0_23_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_16 <= mac_0_23_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_17 <= mac_0_23_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_18 <= mac_0_23_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_19 <= mac_0_23_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_20 <= mac_0_23_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_21 <= mac_0_23_io_mulInput_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_23_io_mulInput_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_23_io_mulInput_sr_22 <= mac_0_23_io_mulInput_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_0 <= io_input_24; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_1 <= mac_0_24_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_2 <= mac_0_24_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_3 <= mac_0_24_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_4 <= mac_0_24_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_5 <= mac_0_24_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_6 <= mac_0_24_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_7 <= mac_0_24_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_8 <= mac_0_24_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_9 <= mac_0_24_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_10 <= mac_0_24_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_11 <= mac_0_24_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_12 <= mac_0_24_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_13 <= mac_0_24_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_14 <= mac_0_24_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_15 <= mac_0_24_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_16 <= mac_0_24_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_17 <= mac_0_24_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_18 <= mac_0_24_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_19 <= mac_0_24_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_20 <= mac_0_24_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_21 <= mac_0_24_io_mulInput_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_22 <= mac_0_24_io_mulInput_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_24_io_mulInput_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_24_io_mulInput_sr_23 <= mac_0_24_io_mulInput_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_0 <= io_input_25; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_1 <= mac_0_25_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_2 <= mac_0_25_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_3 <= mac_0_25_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_4 <= mac_0_25_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_5 <= mac_0_25_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_6 <= mac_0_25_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_7 <= mac_0_25_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_8 <= mac_0_25_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_9 <= mac_0_25_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_10 <= mac_0_25_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_11 <= mac_0_25_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_12 <= mac_0_25_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_13 <= mac_0_25_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_14 <= mac_0_25_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_15 <= mac_0_25_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_16 <= mac_0_25_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_17 <= mac_0_25_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_18 <= mac_0_25_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_19 <= mac_0_25_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_20 <= mac_0_25_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_21 <= mac_0_25_io_mulInput_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_22 <= mac_0_25_io_mulInput_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_23 <= mac_0_25_io_mulInput_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_25_io_mulInput_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_25_io_mulInput_sr_24 <= mac_0_25_io_mulInput_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_0 <= io_input_26; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_1 <= mac_0_26_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_2 <= mac_0_26_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_3 <= mac_0_26_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_4 <= mac_0_26_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_5 <= mac_0_26_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_6 <= mac_0_26_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_7 <= mac_0_26_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_8 <= mac_0_26_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_9 <= mac_0_26_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_10 <= mac_0_26_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_11 <= mac_0_26_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_12 <= mac_0_26_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_13 <= mac_0_26_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_14 <= mac_0_26_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_15 <= mac_0_26_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_16 <= mac_0_26_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_17 <= mac_0_26_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_18 <= mac_0_26_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_19 <= mac_0_26_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_20 <= mac_0_26_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_21 <= mac_0_26_io_mulInput_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_22 <= mac_0_26_io_mulInput_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_23 <= mac_0_26_io_mulInput_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_24 <= mac_0_26_io_mulInput_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_26_io_mulInput_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_26_io_mulInput_sr_25 <= mac_0_26_io_mulInput_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_0 <= io_input_27; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_1 <= mac_0_27_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_2 <= mac_0_27_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_3 <= mac_0_27_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_4 <= mac_0_27_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_5 <= mac_0_27_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_6 <= mac_0_27_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_7 <= mac_0_27_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_8 <= mac_0_27_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_9 <= mac_0_27_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_10 <= mac_0_27_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_11 <= mac_0_27_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_12 <= mac_0_27_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_13 <= mac_0_27_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_14 <= mac_0_27_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_15 <= mac_0_27_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_16 <= mac_0_27_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_17 <= mac_0_27_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_18 <= mac_0_27_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_19 <= mac_0_27_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_20 <= mac_0_27_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_21 <= mac_0_27_io_mulInput_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_22 <= mac_0_27_io_mulInput_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_23 <= mac_0_27_io_mulInput_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_24 <= mac_0_27_io_mulInput_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_25 <= mac_0_27_io_mulInput_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_27_io_mulInput_sr_26 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_27_io_mulInput_sr_26 <= mac_0_27_io_mulInput_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_0 <= io_input_28; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_1 <= mac_0_28_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_2 <= mac_0_28_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_3 <= mac_0_28_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_4 <= mac_0_28_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_5 <= mac_0_28_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_6 <= mac_0_28_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_7 <= mac_0_28_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_8 <= mac_0_28_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_9 <= mac_0_28_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_10 <= mac_0_28_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_11 <= mac_0_28_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_12 <= mac_0_28_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_13 <= mac_0_28_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_14 <= mac_0_28_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_15 <= mac_0_28_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_16 <= mac_0_28_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_17 <= mac_0_28_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_18 <= mac_0_28_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_19 <= mac_0_28_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_20 <= mac_0_28_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_21 <= mac_0_28_io_mulInput_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_22 <= mac_0_28_io_mulInput_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_23 <= mac_0_28_io_mulInput_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_24 <= mac_0_28_io_mulInput_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_25 <= mac_0_28_io_mulInput_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_26 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_26 <= mac_0_28_io_mulInput_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_28_io_mulInput_sr_27 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_28_io_mulInput_sr_27 <= mac_0_28_io_mulInput_sr_26; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_0 <= io_input_29; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_1 <= mac_0_29_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_2 <= mac_0_29_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_3 <= mac_0_29_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_4 <= mac_0_29_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_5 <= mac_0_29_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_6 <= mac_0_29_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_7 <= mac_0_29_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_8 <= mac_0_29_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_9 <= mac_0_29_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_10 <= mac_0_29_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_11 <= mac_0_29_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_12 <= mac_0_29_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_13 <= mac_0_29_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_14 <= mac_0_29_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_15 <= mac_0_29_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_16 <= mac_0_29_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_17 <= mac_0_29_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_18 <= mac_0_29_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_19 <= mac_0_29_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_20 <= mac_0_29_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_21 <= mac_0_29_io_mulInput_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_22 <= mac_0_29_io_mulInput_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_23 <= mac_0_29_io_mulInput_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_24 <= mac_0_29_io_mulInput_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_25 <= mac_0_29_io_mulInput_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_26 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_26 <= mac_0_29_io_mulInput_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_27 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_27 <= mac_0_29_io_mulInput_sr_26; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_29_io_mulInput_sr_28 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_29_io_mulInput_sr_28 <= mac_0_29_io_mulInput_sr_27; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_0 <= io_input_30; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_1 <= mac_0_30_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_2 <= mac_0_30_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_3 <= mac_0_30_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_4 <= mac_0_30_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_5 <= mac_0_30_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_6 <= mac_0_30_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_7 <= mac_0_30_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_8 <= mac_0_30_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_9 <= mac_0_30_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_10 <= mac_0_30_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_11 <= mac_0_30_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_12 <= mac_0_30_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_13 <= mac_0_30_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_14 <= mac_0_30_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_15 <= mac_0_30_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_16 <= mac_0_30_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_17 <= mac_0_30_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_18 <= mac_0_30_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_19 <= mac_0_30_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_20 <= mac_0_30_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_21 <= mac_0_30_io_mulInput_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_22 <= mac_0_30_io_mulInput_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_23 <= mac_0_30_io_mulInput_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_24 <= mac_0_30_io_mulInput_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_25 <= mac_0_30_io_mulInput_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_26 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_26 <= mac_0_30_io_mulInput_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_27 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_27 <= mac_0_30_io_mulInput_sr_26; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_28 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_28 <= mac_0_30_io_mulInput_sr_27; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_30_io_mulInput_sr_29 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_30_io_mulInput_sr_29 <= mac_0_30_io_mulInput_sr_28; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_0 <= io_input_31; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_1 <= mac_0_31_io_mulInput_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_2 <= mac_0_31_io_mulInput_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_3 <= mac_0_31_io_mulInput_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_4 <= mac_0_31_io_mulInput_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_5 <= mac_0_31_io_mulInput_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_6 <= mac_0_31_io_mulInput_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_7 <= mac_0_31_io_mulInput_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_8 <= mac_0_31_io_mulInput_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_9 <= mac_0_31_io_mulInput_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_10 <= mac_0_31_io_mulInput_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_11 <= mac_0_31_io_mulInput_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_12 <= mac_0_31_io_mulInput_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_13 <= mac_0_31_io_mulInput_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_14 <= mac_0_31_io_mulInput_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_15 <= mac_0_31_io_mulInput_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_16 <= mac_0_31_io_mulInput_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_17 <= mac_0_31_io_mulInput_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_18 <= mac_0_31_io_mulInput_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_19 <= mac_0_31_io_mulInput_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_20 <= mac_0_31_io_mulInput_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_21 <= mac_0_31_io_mulInput_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_22 <= mac_0_31_io_mulInput_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_23 <= mac_0_31_io_mulInput_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_24 <= mac_0_31_io_mulInput_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_25 <= mac_0_31_io_mulInput_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_26 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_26 <= mac_0_31_io_mulInput_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_27 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_27 <= mac_0_31_io_mulInput_sr_26; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_28 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_28 <= mac_0_31_io_mulInput_sr_27; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_29 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_29 <= mac_0_31_io_mulInput_sr_28; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      mac_0_31_io_mulInput_sr_30 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      mac_0_31_io_mulInput_sr_30 <= mac_0_31_io_mulInput_sr_29; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_0 <= mac_0_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_1 <= io_output_0_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_2 <= io_output_0_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_3 <= io_output_0_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_4 <= io_output_0_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_5 <= io_output_0_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_6 <= io_output_0_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_7 <= io_output_0_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_8 <= io_output_0_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_9 <= io_output_0_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_10 <= io_output_0_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_11 <= io_output_0_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_12 <= io_output_0_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_13 <= io_output_0_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_14 <= io_output_0_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_15 <= io_output_0_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_16 <= io_output_0_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_17 <= io_output_0_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_18 <= io_output_0_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_19 <= io_output_0_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_20 <= io_output_0_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_21 <= io_output_0_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_22 <= io_output_0_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_23 <= io_output_0_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_24 <= io_output_0_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_25 <= io_output_0_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_26 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_26 <= io_output_0_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_27 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_27 <= io_output_0_sr_26; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_28 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_28 <= io_output_0_sr_27; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_29 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_29 <= io_output_0_sr_28; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_0_sr_30 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_0_sr_30 <= io_output_0_sr_29; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_0 <= mac_1_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_1 <= io_output_1_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_2 <= io_output_1_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_3 <= io_output_1_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_4 <= io_output_1_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_5 <= io_output_1_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_6 <= io_output_1_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_7 <= io_output_1_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_8 <= io_output_1_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_9 <= io_output_1_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_10 <= io_output_1_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_11 <= io_output_1_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_12 <= io_output_1_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_13 <= io_output_1_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_14 <= io_output_1_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_15 <= io_output_1_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_16 <= io_output_1_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_17 <= io_output_1_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_18 <= io_output_1_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_19 <= io_output_1_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_20 <= io_output_1_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_21 <= io_output_1_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_22 <= io_output_1_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_23 <= io_output_1_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_24 <= io_output_1_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_25 <= io_output_1_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_26 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_26 <= io_output_1_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_27 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_27 <= io_output_1_sr_26; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_28 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_28 <= io_output_1_sr_27; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_1_sr_29 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_1_sr_29 <= io_output_1_sr_28; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_0 <= mac_2_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_1 <= io_output_2_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_2 <= io_output_2_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_3 <= io_output_2_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_4 <= io_output_2_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_5 <= io_output_2_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_6 <= io_output_2_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_7 <= io_output_2_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_8 <= io_output_2_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_9 <= io_output_2_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_10 <= io_output_2_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_11 <= io_output_2_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_12 <= io_output_2_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_13 <= io_output_2_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_14 <= io_output_2_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_15 <= io_output_2_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_16 <= io_output_2_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_17 <= io_output_2_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_18 <= io_output_2_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_19 <= io_output_2_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_20 <= io_output_2_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_21 <= io_output_2_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_22 <= io_output_2_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_23 <= io_output_2_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_24 <= io_output_2_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_25 <= io_output_2_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_26 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_26 <= io_output_2_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_27 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_27 <= io_output_2_sr_26; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_2_sr_28 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_2_sr_28 <= io_output_2_sr_27; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_0 <= mac_3_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_1 <= io_output_3_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_2 <= io_output_3_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_3 <= io_output_3_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_4 <= io_output_3_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_5 <= io_output_3_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_6 <= io_output_3_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_7 <= io_output_3_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_8 <= io_output_3_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_9 <= io_output_3_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_10 <= io_output_3_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_11 <= io_output_3_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_12 <= io_output_3_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_13 <= io_output_3_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_14 <= io_output_3_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_15 <= io_output_3_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_16 <= io_output_3_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_17 <= io_output_3_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_18 <= io_output_3_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_19 <= io_output_3_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_20 <= io_output_3_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_21 <= io_output_3_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_22 <= io_output_3_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_23 <= io_output_3_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_24 <= io_output_3_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_25 <= io_output_3_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_26 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_26 <= io_output_3_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_3_sr_27 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_3_sr_27 <= io_output_3_sr_26; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_0 <= mac_4_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_1 <= io_output_4_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_2 <= io_output_4_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_3 <= io_output_4_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_4 <= io_output_4_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_5 <= io_output_4_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_6 <= io_output_4_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_7 <= io_output_4_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_8 <= io_output_4_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_9 <= io_output_4_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_10 <= io_output_4_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_11 <= io_output_4_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_12 <= io_output_4_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_13 <= io_output_4_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_14 <= io_output_4_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_15 <= io_output_4_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_16 <= io_output_4_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_17 <= io_output_4_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_18 <= io_output_4_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_19 <= io_output_4_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_20 <= io_output_4_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_21 <= io_output_4_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_22 <= io_output_4_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_23 <= io_output_4_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_24 <= io_output_4_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_25 <= io_output_4_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_4_sr_26 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_4_sr_26 <= io_output_4_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_0 <= mac_5_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_1 <= io_output_5_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_2 <= io_output_5_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_3 <= io_output_5_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_4 <= io_output_5_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_5 <= io_output_5_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_6 <= io_output_5_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_7 <= io_output_5_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_8 <= io_output_5_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_9 <= io_output_5_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_10 <= io_output_5_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_11 <= io_output_5_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_12 <= io_output_5_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_13 <= io_output_5_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_14 <= io_output_5_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_15 <= io_output_5_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_16 <= io_output_5_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_17 <= io_output_5_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_18 <= io_output_5_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_19 <= io_output_5_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_20 <= io_output_5_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_21 <= io_output_5_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_22 <= io_output_5_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_23 <= io_output_5_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_24 <= io_output_5_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_5_sr_25 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_5_sr_25 <= io_output_5_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_0 <= mac_6_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_1 <= io_output_6_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_2 <= io_output_6_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_3 <= io_output_6_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_4 <= io_output_6_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_5 <= io_output_6_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_6 <= io_output_6_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_7 <= io_output_6_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_8 <= io_output_6_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_9 <= io_output_6_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_10 <= io_output_6_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_11 <= io_output_6_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_12 <= io_output_6_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_13 <= io_output_6_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_14 <= io_output_6_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_15 <= io_output_6_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_16 <= io_output_6_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_17 <= io_output_6_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_18 <= io_output_6_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_19 <= io_output_6_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_20 <= io_output_6_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_21 <= io_output_6_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_22 <= io_output_6_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_23 <= io_output_6_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_6_sr_24 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_6_sr_24 <= io_output_6_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_0 <= mac_7_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_1 <= io_output_7_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_2 <= io_output_7_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_3 <= io_output_7_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_4 <= io_output_7_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_5 <= io_output_7_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_6 <= io_output_7_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_7 <= io_output_7_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_8 <= io_output_7_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_9 <= io_output_7_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_10 <= io_output_7_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_11 <= io_output_7_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_12 <= io_output_7_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_13 <= io_output_7_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_14 <= io_output_7_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_15 <= io_output_7_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_16 <= io_output_7_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_17 <= io_output_7_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_18 <= io_output_7_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_19 <= io_output_7_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_20 <= io_output_7_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_21 <= io_output_7_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_22 <= io_output_7_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_7_sr_23 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_7_sr_23 <= io_output_7_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_0 <= mac_8_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_1 <= io_output_8_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_2 <= io_output_8_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_3 <= io_output_8_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_4 <= io_output_8_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_5 <= io_output_8_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_6 <= io_output_8_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_7 <= io_output_8_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_8 <= io_output_8_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_9 <= io_output_8_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_10 <= io_output_8_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_11 <= io_output_8_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_12 <= io_output_8_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_13 <= io_output_8_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_14 <= io_output_8_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_15 <= io_output_8_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_16 <= io_output_8_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_17 <= io_output_8_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_18 <= io_output_8_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_19 <= io_output_8_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_20 <= io_output_8_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_21 <= io_output_8_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_8_sr_22 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_8_sr_22 <= io_output_8_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_0 <= mac_9_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_1 <= io_output_9_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_2 <= io_output_9_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_3 <= io_output_9_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_4 <= io_output_9_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_5 <= io_output_9_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_6 <= io_output_9_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_7 <= io_output_9_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_8 <= io_output_9_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_9 <= io_output_9_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_10 <= io_output_9_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_11 <= io_output_9_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_12 <= io_output_9_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_13 <= io_output_9_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_14 <= io_output_9_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_15 <= io_output_9_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_16 <= io_output_9_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_17 <= io_output_9_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_18 <= io_output_9_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_19 <= io_output_9_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_20 <= io_output_9_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_9_sr_21 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_9_sr_21 <= io_output_9_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_0 <= mac_10_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_1 <= io_output_10_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_2 <= io_output_10_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_3 <= io_output_10_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_4 <= io_output_10_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_5 <= io_output_10_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_6 <= io_output_10_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_7 <= io_output_10_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_8 <= io_output_10_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_9 <= io_output_10_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_10 <= io_output_10_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_11 <= io_output_10_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_12 <= io_output_10_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_13 <= io_output_10_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_14 <= io_output_10_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_15 <= io_output_10_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_16 <= io_output_10_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_17 <= io_output_10_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_18 <= io_output_10_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_19 <= io_output_10_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_10_sr_20 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_10_sr_20 <= io_output_10_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_0 <= mac_11_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_1 <= io_output_11_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_2 <= io_output_11_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_3 <= io_output_11_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_4 <= io_output_11_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_5 <= io_output_11_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_6 <= io_output_11_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_7 <= io_output_11_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_8 <= io_output_11_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_9 <= io_output_11_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_10 <= io_output_11_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_11 <= io_output_11_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_12 <= io_output_11_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_13 <= io_output_11_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_14 <= io_output_11_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_15 <= io_output_11_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_16 <= io_output_11_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_17 <= io_output_11_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_18 <= io_output_11_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_11_sr_19 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_11_sr_19 <= io_output_11_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_0 <= mac_12_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_1 <= io_output_12_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_2 <= io_output_12_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_3 <= io_output_12_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_4 <= io_output_12_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_5 <= io_output_12_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_6 <= io_output_12_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_7 <= io_output_12_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_8 <= io_output_12_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_9 <= io_output_12_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_10 <= io_output_12_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_11 <= io_output_12_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_12 <= io_output_12_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_13 <= io_output_12_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_14 <= io_output_12_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_15 <= io_output_12_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_16 <= io_output_12_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_17 <= io_output_12_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_12_sr_18 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_12_sr_18 <= io_output_12_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_0 <= mac_13_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_1 <= io_output_13_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_2 <= io_output_13_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_3 <= io_output_13_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_4 <= io_output_13_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_5 <= io_output_13_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_6 <= io_output_13_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_7 <= io_output_13_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_8 <= io_output_13_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_9 <= io_output_13_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_10 <= io_output_13_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_11 <= io_output_13_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_12 <= io_output_13_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_13 <= io_output_13_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_14 <= io_output_13_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_15 <= io_output_13_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_16 <= io_output_13_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_13_sr_17 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_13_sr_17 <= io_output_13_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_0 <= mac_14_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_1 <= io_output_14_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_2 <= io_output_14_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_3 <= io_output_14_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_4 <= io_output_14_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_5 <= io_output_14_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_6 <= io_output_14_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_7 <= io_output_14_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_8 <= io_output_14_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_9 <= io_output_14_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_10 <= io_output_14_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_11 <= io_output_14_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_12 <= io_output_14_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_13 <= io_output_14_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_14 <= io_output_14_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_15 <= io_output_14_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_14_sr_16 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_14_sr_16 <= io_output_14_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_0 <= mac_15_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_1 <= io_output_15_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_2 <= io_output_15_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_3 <= io_output_15_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_4 <= io_output_15_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_5 <= io_output_15_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_6 <= io_output_15_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_7 <= io_output_15_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_8 <= io_output_15_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_9 <= io_output_15_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_10 <= io_output_15_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_11 <= io_output_15_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_12 <= io_output_15_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_13 <= io_output_15_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_14 <= io_output_15_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_15_sr_15 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_15_sr_15 <= io_output_15_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_0 <= mac_16_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_1 <= io_output_16_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_2 <= io_output_16_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_3 <= io_output_16_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_4 <= io_output_16_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_5 <= io_output_16_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_6 <= io_output_16_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_7 <= io_output_16_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_8 <= io_output_16_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_9 <= io_output_16_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_10 <= io_output_16_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_11 <= io_output_16_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_12 <= io_output_16_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_13 <= io_output_16_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_16_sr_14 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_16_sr_14 <= io_output_16_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_0 <= mac_17_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_1 <= io_output_17_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_2 <= io_output_17_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_3 <= io_output_17_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_4 <= io_output_17_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_5 <= io_output_17_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_6 <= io_output_17_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_7 <= io_output_17_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_8 <= io_output_17_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_9 <= io_output_17_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_10 <= io_output_17_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_11 <= io_output_17_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_12 <= io_output_17_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_17_sr_13 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_17_sr_13 <= io_output_17_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_0 <= mac_18_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_1 <= io_output_18_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_2 <= io_output_18_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_3 <= io_output_18_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_4 <= io_output_18_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_5 <= io_output_18_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_6 <= io_output_18_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_7 <= io_output_18_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_8 <= io_output_18_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_9 <= io_output_18_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_10 <= io_output_18_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_11 <= io_output_18_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_18_sr_12 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_18_sr_12 <= io_output_18_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_0 <= mac_19_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_1 <= io_output_19_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_2 <= io_output_19_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_3 <= io_output_19_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_4 <= io_output_19_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_5 <= io_output_19_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_6 <= io_output_19_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_7 <= io_output_19_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_8 <= io_output_19_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_9 <= io_output_19_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_10 <= io_output_19_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_19_sr_11 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_19_sr_11 <= io_output_19_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_0 <= mac_20_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_1 <= io_output_20_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_2 <= io_output_20_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_3 <= io_output_20_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_4 <= io_output_20_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_5 <= io_output_20_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_6 <= io_output_20_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_7 <= io_output_20_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_8 <= io_output_20_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_9 <= io_output_20_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_20_sr_10 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_20_sr_10 <= io_output_20_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_21_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_21_sr_0 <= mac_21_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_21_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_21_sr_1 <= io_output_21_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_21_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_21_sr_2 <= io_output_21_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_21_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_21_sr_3 <= io_output_21_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_21_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_21_sr_4 <= io_output_21_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_21_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_21_sr_5 <= io_output_21_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_21_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_21_sr_6 <= io_output_21_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_21_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_21_sr_7 <= io_output_21_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_21_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_21_sr_8 <= io_output_21_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_21_sr_9 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_21_sr_9 <= io_output_21_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_22_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_22_sr_0 <= mac_22_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_22_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_22_sr_1 <= io_output_22_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_22_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_22_sr_2 <= io_output_22_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_22_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_22_sr_3 <= io_output_22_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_22_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_22_sr_4 <= io_output_22_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_22_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_22_sr_5 <= io_output_22_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_22_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_22_sr_6 <= io_output_22_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_22_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_22_sr_7 <= io_output_22_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_22_sr_8 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_22_sr_8 <= io_output_22_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_23_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_23_sr_0 <= mac_23_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_23_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_23_sr_1 <= io_output_23_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_23_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_23_sr_2 <= io_output_23_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_23_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_23_sr_3 <= io_output_23_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_23_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_23_sr_4 <= io_output_23_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_23_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_23_sr_5 <= io_output_23_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_23_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_23_sr_6 <= io_output_23_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_23_sr_7 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_23_sr_7 <= io_output_23_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_24_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_24_sr_0 <= mac_24_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_24_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_24_sr_1 <= io_output_24_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_24_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_24_sr_2 <= io_output_24_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_24_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_24_sr_3 <= io_output_24_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_24_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_24_sr_4 <= io_output_24_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_24_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_24_sr_5 <= io_output_24_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_24_sr_6 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_24_sr_6 <= io_output_24_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_25_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_25_sr_0 <= mac_25_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_25_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_25_sr_1 <= io_output_25_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_25_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_25_sr_2 <= io_output_25_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_25_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_25_sr_3 <= io_output_25_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_25_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_25_sr_4 <= io_output_25_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_25_sr_5 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_25_sr_5 <= io_output_25_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_26_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_26_sr_0 <= mac_26_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_26_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_26_sr_1 <= io_output_26_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_26_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_26_sr_2 <= io_output_26_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_26_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_26_sr_3 <= io_output_26_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_26_sr_4 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_26_sr_4 <= io_output_26_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_27_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_27_sr_0 <= mac_27_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_27_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_27_sr_1 <= io_output_27_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_27_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_27_sr_2 <= io_output_27_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_27_sr_3 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_27_sr_3 <= io_output_27_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_28_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_28_sr_0 <= mac_28_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_28_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_28_sr_1 <= io_output_28_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_28_sr_2 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_28_sr_2 <= io_output_28_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_29_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_29_sr_0 <= mac_29_31_io_output; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_29_sr_1 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_29_sr_1 <= io_output_29_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      io_output_30_sr_0 <= 16'sh0; // @[ShiftRegister.scala 10:22]
    end else begin
      io_output_30_sr_0 <= mac_30_31_io_output; // @[ShiftRegister.scala 25:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bias_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  bias_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  bias_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  bias_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  bias_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  bias_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  bias_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  bias_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  bias_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  bias_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  bias_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  bias_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  bias_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  bias_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  bias_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  bias_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  bias_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  bias_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  bias_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  bias_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  bias_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  bias_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  bias_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  bias_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  bias_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  bias_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  bias_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  bias_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  bias_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  bias_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  bias_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  bias_31 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  mac_0_1_io_mulInput_sr_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  mac_0_2_io_mulInput_sr_0 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  mac_0_2_io_mulInput_sr_1 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  mac_0_3_io_mulInput_sr_0 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  mac_0_3_io_mulInput_sr_1 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  mac_0_3_io_mulInput_sr_2 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  mac_0_4_io_mulInput_sr_0 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  mac_0_4_io_mulInput_sr_1 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  mac_0_4_io_mulInput_sr_2 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  mac_0_4_io_mulInput_sr_3 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  mac_0_5_io_mulInput_sr_0 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  mac_0_5_io_mulInput_sr_1 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  mac_0_5_io_mulInput_sr_2 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  mac_0_5_io_mulInput_sr_3 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  mac_0_5_io_mulInput_sr_4 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  mac_0_6_io_mulInput_sr_0 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  mac_0_6_io_mulInput_sr_1 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  mac_0_6_io_mulInput_sr_2 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  mac_0_6_io_mulInput_sr_3 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  mac_0_6_io_mulInput_sr_4 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  mac_0_6_io_mulInput_sr_5 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  mac_0_7_io_mulInput_sr_0 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  mac_0_7_io_mulInput_sr_1 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  mac_0_7_io_mulInput_sr_2 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  mac_0_7_io_mulInput_sr_3 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  mac_0_7_io_mulInput_sr_4 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  mac_0_7_io_mulInput_sr_5 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  mac_0_7_io_mulInput_sr_6 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  mac_0_8_io_mulInput_sr_0 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  mac_0_8_io_mulInput_sr_1 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  mac_0_8_io_mulInput_sr_2 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  mac_0_8_io_mulInput_sr_3 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  mac_0_8_io_mulInput_sr_4 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  mac_0_8_io_mulInput_sr_5 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  mac_0_8_io_mulInput_sr_6 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  mac_0_8_io_mulInput_sr_7 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  mac_0_9_io_mulInput_sr_0 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  mac_0_9_io_mulInput_sr_1 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  mac_0_9_io_mulInput_sr_2 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  mac_0_9_io_mulInput_sr_3 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  mac_0_9_io_mulInput_sr_4 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  mac_0_9_io_mulInput_sr_5 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  mac_0_9_io_mulInput_sr_6 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  mac_0_9_io_mulInput_sr_7 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  mac_0_9_io_mulInput_sr_8 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  mac_0_10_io_mulInput_sr_0 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  mac_0_10_io_mulInput_sr_1 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  mac_0_10_io_mulInput_sr_2 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  mac_0_10_io_mulInput_sr_3 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  mac_0_10_io_mulInput_sr_4 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  mac_0_10_io_mulInput_sr_5 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  mac_0_10_io_mulInput_sr_6 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  mac_0_10_io_mulInput_sr_7 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  mac_0_10_io_mulInput_sr_8 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  mac_0_10_io_mulInput_sr_9 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_0 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_1 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_2 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_3 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_4 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_5 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_6 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_7 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_8 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_9 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  mac_0_11_io_mulInput_sr_10 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_0 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_1 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_2 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_3 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_4 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_5 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_6 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_7 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_8 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_9 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_10 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  mac_0_12_io_mulInput_sr_11 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_0 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_1 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_2 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_3 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_4 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_5 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_6 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_7 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_8 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_9 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_10 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_11 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  mac_0_13_io_mulInput_sr_12 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_0 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_1 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_2 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_3 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_4 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_5 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_6 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_7 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_8 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_9 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_10 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_11 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_12 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  mac_0_14_io_mulInput_sr_13 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_0 = _RAND_137[15:0];
  _RAND_138 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_1 = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_2 = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_3 = _RAND_140[15:0];
  _RAND_141 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_4 = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_5 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_6 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_7 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_8 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_9 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_10 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_11 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_12 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_13 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  mac_0_15_io_mulInput_sr_14 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_0 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_1 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_2 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_3 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_4 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_5 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_6 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_7 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_8 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_9 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_10 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_11 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_12 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_13 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_14 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  mac_0_16_io_mulInput_sr_15 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_0 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_1 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_2 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_3 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_4 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_5 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_6 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_7 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_8 = _RAND_176[15:0];
  _RAND_177 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_9 = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_10 = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_11 = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_12 = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_13 = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_14 = _RAND_182[15:0];
  _RAND_183 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_15 = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  mac_0_17_io_mulInput_sr_16 = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_0 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_1 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_2 = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_3 = _RAND_188[15:0];
  _RAND_189 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_4 = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_5 = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_6 = _RAND_191[15:0];
  _RAND_192 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_7 = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_8 = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_9 = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_10 = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_11 = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_12 = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_13 = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_14 = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_15 = _RAND_200[15:0];
  _RAND_201 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_16 = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  mac_0_18_io_mulInput_sr_17 = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_0 = _RAND_203[15:0];
  _RAND_204 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_1 = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_2 = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_3 = _RAND_206[15:0];
  _RAND_207 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_4 = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_5 = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_6 = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_7 = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_8 = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_9 = _RAND_212[15:0];
  _RAND_213 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_10 = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_11 = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_12 = _RAND_215[15:0];
  _RAND_216 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_13 = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_14 = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_15 = _RAND_218[15:0];
  _RAND_219 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_16 = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_17 = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  mac_0_19_io_mulInput_sr_18 = _RAND_221[15:0];
  _RAND_222 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_0 = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_1 = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_2 = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_3 = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_4 = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_5 = _RAND_227[15:0];
  _RAND_228 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_6 = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_7 = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_8 = _RAND_230[15:0];
  _RAND_231 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_9 = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_10 = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_11 = _RAND_233[15:0];
  _RAND_234 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_12 = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_13 = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_14 = _RAND_236[15:0];
  _RAND_237 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_15 = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_16 = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_17 = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_18 = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  mac_0_20_io_mulInput_sr_19 = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_0 = _RAND_242[15:0];
  _RAND_243 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_1 = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_2 = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_3 = _RAND_245[15:0];
  _RAND_246 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_4 = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_5 = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_6 = _RAND_248[15:0];
  _RAND_249 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_7 = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_8 = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_9 = _RAND_251[15:0];
  _RAND_252 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_10 = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_11 = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_12 = _RAND_254[15:0];
  _RAND_255 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_13 = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_14 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_15 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_16 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_17 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_18 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_19 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  mac_0_21_io_mulInput_sr_20 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_0 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_1 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_2 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_3 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_4 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_5 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_6 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_7 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_8 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_9 = _RAND_272[15:0];
  _RAND_273 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_10 = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_11 = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_12 = _RAND_275[15:0];
  _RAND_276 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_13 = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_14 = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_15 = _RAND_278[15:0];
  _RAND_279 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_16 = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_17 = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_18 = _RAND_281[15:0];
  _RAND_282 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_19 = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_20 = _RAND_283[15:0];
  _RAND_284 = {1{`RANDOM}};
  mac_0_22_io_mulInput_sr_21 = _RAND_284[15:0];
  _RAND_285 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_0 = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_1 = _RAND_286[15:0];
  _RAND_287 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_2 = _RAND_287[15:0];
  _RAND_288 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_3 = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_4 = _RAND_289[15:0];
  _RAND_290 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_5 = _RAND_290[15:0];
  _RAND_291 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_6 = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_7 = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_8 = _RAND_293[15:0];
  _RAND_294 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_9 = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_10 = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_11 = _RAND_296[15:0];
  _RAND_297 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_12 = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_13 = _RAND_298[15:0];
  _RAND_299 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_14 = _RAND_299[15:0];
  _RAND_300 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_15 = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_16 = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_17 = _RAND_302[15:0];
  _RAND_303 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_18 = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_19 = _RAND_304[15:0];
  _RAND_305 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_20 = _RAND_305[15:0];
  _RAND_306 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_21 = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  mac_0_23_io_mulInput_sr_22 = _RAND_307[15:0];
  _RAND_308 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_0 = _RAND_308[15:0];
  _RAND_309 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_1 = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_2 = _RAND_310[15:0];
  _RAND_311 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_3 = _RAND_311[15:0];
  _RAND_312 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_4 = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_5 = _RAND_313[15:0];
  _RAND_314 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_6 = _RAND_314[15:0];
  _RAND_315 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_7 = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_8 = _RAND_316[15:0];
  _RAND_317 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_9 = _RAND_317[15:0];
  _RAND_318 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_10 = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_11 = _RAND_319[15:0];
  _RAND_320 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_12 = _RAND_320[15:0];
  _RAND_321 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_13 = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_14 = _RAND_322[15:0];
  _RAND_323 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_15 = _RAND_323[15:0];
  _RAND_324 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_16 = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_17 = _RAND_325[15:0];
  _RAND_326 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_18 = _RAND_326[15:0];
  _RAND_327 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_19 = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_20 = _RAND_328[15:0];
  _RAND_329 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_21 = _RAND_329[15:0];
  _RAND_330 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_22 = _RAND_330[15:0];
  _RAND_331 = {1{`RANDOM}};
  mac_0_24_io_mulInput_sr_23 = _RAND_331[15:0];
  _RAND_332 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_0 = _RAND_332[15:0];
  _RAND_333 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_1 = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_2 = _RAND_334[15:0];
  _RAND_335 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_3 = _RAND_335[15:0];
  _RAND_336 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_4 = _RAND_336[15:0];
  _RAND_337 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_5 = _RAND_337[15:0];
  _RAND_338 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_6 = _RAND_338[15:0];
  _RAND_339 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_7 = _RAND_339[15:0];
  _RAND_340 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_8 = _RAND_340[15:0];
  _RAND_341 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_9 = _RAND_341[15:0];
  _RAND_342 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_10 = _RAND_342[15:0];
  _RAND_343 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_11 = _RAND_343[15:0];
  _RAND_344 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_12 = _RAND_344[15:0];
  _RAND_345 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_13 = _RAND_345[15:0];
  _RAND_346 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_14 = _RAND_346[15:0];
  _RAND_347 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_15 = _RAND_347[15:0];
  _RAND_348 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_16 = _RAND_348[15:0];
  _RAND_349 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_17 = _RAND_349[15:0];
  _RAND_350 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_18 = _RAND_350[15:0];
  _RAND_351 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_19 = _RAND_351[15:0];
  _RAND_352 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_20 = _RAND_352[15:0];
  _RAND_353 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_21 = _RAND_353[15:0];
  _RAND_354 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_22 = _RAND_354[15:0];
  _RAND_355 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_23 = _RAND_355[15:0];
  _RAND_356 = {1{`RANDOM}};
  mac_0_25_io_mulInput_sr_24 = _RAND_356[15:0];
  _RAND_357 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_0 = _RAND_357[15:0];
  _RAND_358 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_1 = _RAND_358[15:0];
  _RAND_359 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_2 = _RAND_359[15:0];
  _RAND_360 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_3 = _RAND_360[15:0];
  _RAND_361 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_4 = _RAND_361[15:0];
  _RAND_362 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_5 = _RAND_362[15:0];
  _RAND_363 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_6 = _RAND_363[15:0];
  _RAND_364 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_7 = _RAND_364[15:0];
  _RAND_365 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_8 = _RAND_365[15:0];
  _RAND_366 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_9 = _RAND_366[15:0];
  _RAND_367 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_10 = _RAND_367[15:0];
  _RAND_368 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_11 = _RAND_368[15:0];
  _RAND_369 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_12 = _RAND_369[15:0];
  _RAND_370 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_13 = _RAND_370[15:0];
  _RAND_371 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_14 = _RAND_371[15:0];
  _RAND_372 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_15 = _RAND_372[15:0];
  _RAND_373 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_16 = _RAND_373[15:0];
  _RAND_374 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_17 = _RAND_374[15:0];
  _RAND_375 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_18 = _RAND_375[15:0];
  _RAND_376 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_19 = _RAND_376[15:0];
  _RAND_377 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_20 = _RAND_377[15:0];
  _RAND_378 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_21 = _RAND_378[15:0];
  _RAND_379 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_22 = _RAND_379[15:0];
  _RAND_380 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_23 = _RAND_380[15:0];
  _RAND_381 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_24 = _RAND_381[15:0];
  _RAND_382 = {1{`RANDOM}};
  mac_0_26_io_mulInput_sr_25 = _RAND_382[15:0];
  _RAND_383 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_0 = _RAND_383[15:0];
  _RAND_384 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_1 = _RAND_384[15:0];
  _RAND_385 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_2 = _RAND_385[15:0];
  _RAND_386 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_3 = _RAND_386[15:0];
  _RAND_387 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_4 = _RAND_387[15:0];
  _RAND_388 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_5 = _RAND_388[15:0];
  _RAND_389 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_6 = _RAND_389[15:0];
  _RAND_390 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_7 = _RAND_390[15:0];
  _RAND_391 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_8 = _RAND_391[15:0];
  _RAND_392 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_9 = _RAND_392[15:0];
  _RAND_393 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_10 = _RAND_393[15:0];
  _RAND_394 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_11 = _RAND_394[15:0];
  _RAND_395 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_12 = _RAND_395[15:0];
  _RAND_396 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_13 = _RAND_396[15:0];
  _RAND_397 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_14 = _RAND_397[15:0];
  _RAND_398 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_15 = _RAND_398[15:0];
  _RAND_399 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_16 = _RAND_399[15:0];
  _RAND_400 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_17 = _RAND_400[15:0];
  _RAND_401 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_18 = _RAND_401[15:0];
  _RAND_402 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_19 = _RAND_402[15:0];
  _RAND_403 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_20 = _RAND_403[15:0];
  _RAND_404 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_21 = _RAND_404[15:0];
  _RAND_405 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_22 = _RAND_405[15:0];
  _RAND_406 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_23 = _RAND_406[15:0];
  _RAND_407 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_24 = _RAND_407[15:0];
  _RAND_408 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_25 = _RAND_408[15:0];
  _RAND_409 = {1{`RANDOM}};
  mac_0_27_io_mulInput_sr_26 = _RAND_409[15:0];
  _RAND_410 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_0 = _RAND_410[15:0];
  _RAND_411 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_1 = _RAND_411[15:0];
  _RAND_412 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_2 = _RAND_412[15:0];
  _RAND_413 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_3 = _RAND_413[15:0];
  _RAND_414 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_4 = _RAND_414[15:0];
  _RAND_415 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_5 = _RAND_415[15:0];
  _RAND_416 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_6 = _RAND_416[15:0];
  _RAND_417 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_7 = _RAND_417[15:0];
  _RAND_418 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_8 = _RAND_418[15:0];
  _RAND_419 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_9 = _RAND_419[15:0];
  _RAND_420 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_10 = _RAND_420[15:0];
  _RAND_421 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_11 = _RAND_421[15:0];
  _RAND_422 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_12 = _RAND_422[15:0];
  _RAND_423 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_13 = _RAND_423[15:0];
  _RAND_424 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_14 = _RAND_424[15:0];
  _RAND_425 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_15 = _RAND_425[15:0];
  _RAND_426 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_16 = _RAND_426[15:0];
  _RAND_427 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_17 = _RAND_427[15:0];
  _RAND_428 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_18 = _RAND_428[15:0];
  _RAND_429 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_19 = _RAND_429[15:0];
  _RAND_430 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_20 = _RAND_430[15:0];
  _RAND_431 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_21 = _RAND_431[15:0];
  _RAND_432 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_22 = _RAND_432[15:0];
  _RAND_433 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_23 = _RAND_433[15:0];
  _RAND_434 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_24 = _RAND_434[15:0];
  _RAND_435 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_25 = _RAND_435[15:0];
  _RAND_436 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_26 = _RAND_436[15:0];
  _RAND_437 = {1{`RANDOM}};
  mac_0_28_io_mulInput_sr_27 = _RAND_437[15:0];
  _RAND_438 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_0 = _RAND_438[15:0];
  _RAND_439 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_1 = _RAND_439[15:0];
  _RAND_440 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_2 = _RAND_440[15:0];
  _RAND_441 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_3 = _RAND_441[15:0];
  _RAND_442 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_4 = _RAND_442[15:0];
  _RAND_443 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_5 = _RAND_443[15:0];
  _RAND_444 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_6 = _RAND_444[15:0];
  _RAND_445 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_7 = _RAND_445[15:0];
  _RAND_446 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_8 = _RAND_446[15:0];
  _RAND_447 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_9 = _RAND_447[15:0];
  _RAND_448 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_10 = _RAND_448[15:0];
  _RAND_449 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_11 = _RAND_449[15:0];
  _RAND_450 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_12 = _RAND_450[15:0];
  _RAND_451 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_13 = _RAND_451[15:0];
  _RAND_452 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_14 = _RAND_452[15:0];
  _RAND_453 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_15 = _RAND_453[15:0];
  _RAND_454 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_16 = _RAND_454[15:0];
  _RAND_455 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_17 = _RAND_455[15:0];
  _RAND_456 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_18 = _RAND_456[15:0];
  _RAND_457 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_19 = _RAND_457[15:0];
  _RAND_458 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_20 = _RAND_458[15:0];
  _RAND_459 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_21 = _RAND_459[15:0];
  _RAND_460 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_22 = _RAND_460[15:0];
  _RAND_461 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_23 = _RAND_461[15:0];
  _RAND_462 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_24 = _RAND_462[15:0];
  _RAND_463 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_25 = _RAND_463[15:0];
  _RAND_464 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_26 = _RAND_464[15:0];
  _RAND_465 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_27 = _RAND_465[15:0];
  _RAND_466 = {1{`RANDOM}};
  mac_0_29_io_mulInput_sr_28 = _RAND_466[15:0];
  _RAND_467 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_0 = _RAND_467[15:0];
  _RAND_468 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_1 = _RAND_468[15:0];
  _RAND_469 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_2 = _RAND_469[15:0];
  _RAND_470 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_3 = _RAND_470[15:0];
  _RAND_471 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_4 = _RAND_471[15:0];
  _RAND_472 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_5 = _RAND_472[15:0];
  _RAND_473 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_6 = _RAND_473[15:0];
  _RAND_474 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_7 = _RAND_474[15:0];
  _RAND_475 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_8 = _RAND_475[15:0];
  _RAND_476 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_9 = _RAND_476[15:0];
  _RAND_477 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_10 = _RAND_477[15:0];
  _RAND_478 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_11 = _RAND_478[15:0];
  _RAND_479 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_12 = _RAND_479[15:0];
  _RAND_480 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_13 = _RAND_480[15:0];
  _RAND_481 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_14 = _RAND_481[15:0];
  _RAND_482 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_15 = _RAND_482[15:0];
  _RAND_483 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_16 = _RAND_483[15:0];
  _RAND_484 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_17 = _RAND_484[15:0];
  _RAND_485 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_18 = _RAND_485[15:0];
  _RAND_486 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_19 = _RAND_486[15:0];
  _RAND_487 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_20 = _RAND_487[15:0];
  _RAND_488 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_21 = _RAND_488[15:0];
  _RAND_489 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_22 = _RAND_489[15:0];
  _RAND_490 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_23 = _RAND_490[15:0];
  _RAND_491 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_24 = _RAND_491[15:0];
  _RAND_492 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_25 = _RAND_492[15:0];
  _RAND_493 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_26 = _RAND_493[15:0];
  _RAND_494 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_27 = _RAND_494[15:0];
  _RAND_495 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_28 = _RAND_495[15:0];
  _RAND_496 = {1{`RANDOM}};
  mac_0_30_io_mulInput_sr_29 = _RAND_496[15:0];
  _RAND_497 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_0 = _RAND_497[15:0];
  _RAND_498 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_1 = _RAND_498[15:0];
  _RAND_499 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_2 = _RAND_499[15:0];
  _RAND_500 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_3 = _RAND_500[15:0];
  _RAND_501 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_4 = _RAND_501[15:0];
  _RAND_502 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_5 = _RAND_502[15:0];
  _RAND_503 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_6 = _RAND_503[15:0];
  _RAND_504 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_7 = _RAND_504[15:0];
  _RAND_505 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_8 = _RAND_505[15:0];
  _RAND_506 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_9 = _RAND_506[15:0];
  _RAND_507 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_10 = _RAND_507[15:0];
  _RAND_508 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_11 = _RAND_508[15:0];
  _RAND_509 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_12 = _RAND_509[15:0];
  _RAND_510 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_13 = _RAND_510[15:0];
  _RAND_511 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_14 = _RAND_511[15:0];
  _RAND_512 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_15 = _RAND_512[15:0];
  _RAND_513 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_16 = _RAND_513[15:0];
  _RAND_514 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_17 = _RAND_514[15:0];
  _RAND_515 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_18 = _RAND_515[15:0];
  _RAND_516 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_19 = _RAND_516[15:0];
  _RAND_517 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_20 = _RAND_517[15:0];
  _RAND_518 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_21 = _RAND_518[15:0];
  _RAND_519 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_22 = _RAND_519[15:0];
  _RAND_520 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_23 = _RAND_520[15:0];
  _RAND_521 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_24 = _RAND_521[15:0];
  _RAND_522 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_25 = _RAND_522[15:0];
  _RAND_523 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_26 = _RAND_523[15:0];
  _RAND_524 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_27 = _RAND_524[15:0];
  _RAND_525 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_28 = _RAND_525[15:0];
  _RAND_526 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_29 = _RAND_526[15:0];
  _RAND_527 = {1{`RANDOM}};
  mac_0_31_io_mulInput_sr_30 = _RAND_527[15:0];
  _RAND_528 = {1{`RANDOM}};
  io_output_0_sr_0 = _RAND_528[15:0];
  _RAND_529 = {1{`RANDOM}};
  io_output_0_sr_1 = _RAND_529[15:0];
  _RAND_530 = {1{`RANDOM}};
  io_output_0_sr_2 = _RAND_530[15:0];
  _RAND_531 = {1{`RANDOM}};
  io_output_0_sr_3 = _RAND_531[15:0];
  _RAND_532 = {1{`RANDOM}};
  io_output_0_sr_4 = _RAND_532[15:0];
  _RAND_533 = {1{`RANDOM}};
  io_output_0_sr_5 = _RAND_533[15:0];
  _RAND_534 = {1{`RANDOM}};
  io_output_0_sr_6 = _RAND_534[15:0];
  _RAND_535 = {1{`RANDOM}};
  io_output_0_sr_7 = _RAND_535[15:0];
  _RAND_536 = {1{`RANDOM}};
  io_output_0_sr_8 = _RAND_536[15:0];
  _RAND_537 = {1{`RANDOM}};
  io_output_0_sr_9 = _RAND_537[15:0];
  _RAND_538 = {1{`RANDOM}};
  io_output_0_sr_10 = _RAND_538[15:0];
  _RAND_539 = {1{`RANDOM}};
  io_output_0_sr_11 = _RAND_539[15:0];
  _RAND_540 = {1{`RANDOM}};
  io_output_0_sr_12 = _RAND_540[15:0];
  _RAND_541 = {1{`RANDOM}};
  io_output_0_sr_13 = _RAND_541[15:0];
  _RAND_542 = {1{`RANDOM}};
  io_output_0_sr_14 = _RAND_542[15:0];
  _RAND_543 = {1{`RANDOM}};
  io_output_0_sr_15 = _RAND_543[15:0];
  _RAND_544 = {1{`RANDOM}};
  io_output_0_sr_16 = _RAND_544[15:0];
  _RAND_545 = {1{`RANDOM}};
  io_output_0_sr_17 = _RAND_545[15:0];
  _RAND_546 = {1{`RANDOM}};
  io_output_0_sr_18 = _RAND_546[15:0];
  _RAND_547 = {1{`RANDOM}};
  io_output_0_sr_19 = _RAND_547[15:0];
  _RAND_548 = {1{`RANDOM}};
  io_output_0_sr_20 = _RAND_548[15:0];
  _RAND_549 = {1{`RANDOM}};
  io_output_0_sr_21 = _RAND_549[15:0];
  _RAND_550 = {1{`RANDOM}};
  io_output_0_sr_22 = _RAND_550[15:0];
  _RAND_551 = {1{`RANDOM}};
  io_output_0_sr_23 = _RAND_551[15:0];
  _RAND_552 = {1{`RANDOM}};
  io_output_0_sr_24 = _RAND_552[15:0];
  _RAND_553 = {1{`RANDOM}};
  io_output_0_sr_25 = _RAND_553[15:0];
  _RAND_554 = {1{`RANDOM}};
  io_output_0_sr_26 = _RAND_554[15:0];
  _RAND_555 = {1{`RANDOM}};
  io_output_0_sr_27 = _RAND_555[15:0];
  _RAND_556 = {1{`RANDOM}};
  io_output_0_sr_28 = _RAND_556[15:0];
  _RAND_557 = {1{`RANDOM}};
  io_output_0_sr_29 = _RAND_557[15:0];
  _RAND_558 = {1{`RANDOM}};
  io_output_0_sr_30 = _RAND_558[15:0];
  _RAND_559 = {1{`RANDOM}};
  io_output_1_sr_0 = _RAND_559[15:0];
  _RAND_560 = {1{`RANDOM}};
  io_output_1_sr_1 = _RAND_560[15:0];
  _RAND_561 = {1{`RANDOM}};
  io_output_1_sr_2 = _RAND_561[15:0];
  _RAND_562 = {1{`RANDOM}};
  io_output_1_sr_3 = _RAND_562[15:0];
  _RAND_563 = {1{`RANDOM}};
  io_output_1_sr_4 = _RAND_563[15:0];
  _RAND_564 = {1{`RANDOM}};
  io_output_1_sr_5 = _RAND_564[15:0];
  _RAND_565 = {1{`RANDOM}};
  io_output_1_sr_6 = _RAND_565[15:0];
  _RAND_566 = {1{`RANDOM}};
  io_output_1_sr_7 = _RAND_566[15:0];
  _RAND_567 = {1{`RANDOM}};
  io_output_1_sr_8 = _RAND_567[15:0];
  _RAND_568 = {1{`RANDOM}};
  io_output_1_sr_9 = _RAND_568[15:0];
  _RAND_569 = {1{`RANDOM}};
  io_output_1_sr_10 = _RAND_569[15:0];
  _RAND_570 = {1{`RANDOM}};
  io_output_1_sr_11 = _RAND_570[15:0];
  _RAND_571 = {1{`RANDOM}};
  io_output_1_sr_12 = _RAND_571[15:0];
  _RAND_572 = {1{`RANDOM}};
  io_output_1_sr_13 = _RAND_572[15:0];
  _RAND_573 = {1{`RANDOM}};
  io_output_1_sr_14 = _RAND_573[15:0];
  _RAND_574 = {1{`RANDOM}};
  io_output_1_sr_15 = _RAND_574[15:0];
  _RAND_575 = {1{`RANDOM}};
  io_output_1_sr_16 = _RAND_575[15:0];
  _RAND_576 = {1{`RANDOM}};
  io_output_1_sr_17 = _RAND_576[15:0];
  _RAND_577 = {1{`RANDOM}};
  io_output_1_sr_18 = _RAND_577[15:0];
  _RAND_578 = {1{`RANDOM}};
  io_output_1_sr_19 = _RAND_578[15:0];
  _RAND_579 = {1{`RANDOM}};
  io_output_1_sr_20 = _RAND_579[15:0];
  _RAND_580 = {1{`RANDOM}};
  io_output_1_sr_21 = _RAND_580[15:0];
  _RAND_581 = {1{`RANDOM}};
  io_output_1_sr_22 = _RAND_581[15:0];
  _RAND_582 = {1{`RANDOM}};
  io_output_1_sr_23 = _RAND_582[15:0];
  _RAND_583 = {1{`RANDOM}};
  io_output_1_sr_24 = _RAND_583[15:0];
  _RAND_584 = {1{`RANDOM}};
  io_output_1_sr_25 = _RAND_584[15:0];
  _RAND_585 = {1{`RANDOM}};
  io_output_1_sr_26 = _RAND_585[15:0];
  _RAND_586 = {1{`RANDOM}};
  io_output_1_sr_27 = _RAND_586[15:0];
  _RAND_587 = {1{`RANDOM}};
  io_output_1_sr_28 = _RAND_587[15:0];
  _RAND_588 = {1{`RANDOM}};
  io_output_1_sr_29 = _RAND_588[15:0];
  _RAND_589 = {1{`RANDOM}};
  io_output_2_sr_0 = _RAND_589[15:0];
  _RAND_590 = {1{`RANDOM}};
  io_output_2_sr_1 = _RAND_590[15:0];
  _RAND_591 = {1{`RANDOM}};
  io_output_2_sr_2 = _RAND_591[15:0];
  _RAND_592 = {1{`RANDOM}};
  io_output_2_sr_3 = _RAND_592[15:0];
  _RAND_593 = {1{`RANDOM}};
  io_output_2_sr_4 = _RAND_593[15:0];
  _RAND_594 = {1{`RANDOM}};
  io_output_2_sr_5 = _RAND_594[15:0];
  _RAND_595 = {1{`RANDOM}};
  io_output_2_sr_6 = _RAND_595[15:0];
  _RAND_596 = {1{`RANDOM}};
  io_output_2_sr_7 = _RAND_596[15:0];
  _RAND_597 = {1{`RANDOM}};
  io_output_2_sr_8 = _RAND_597[15:0];
  _RAND_598 = {1{`RANDOM}};
  io_output_2_sr_9 = _RAND_598[15:0];
  _RAND_599 = {1{`RANDOM}};
  io_output_2_sr_10 = _RAND_599[15:0];
  _RAND_600 = {1{`RANDOM}};
  io_output_2_sr_11 = _RAND_600[15:0];
  _RAND_601 = {1{`RANDOM}};
  io_output_2_sr_12 = _RAND_601[15:0];
  _RAND_602 = {1{`RANDOM}};
  io_output_2_sr_13 = _RAND_602[15:0];
  _RAND_603 = {1{`RANDOM}};
  io_output_2_sr_14 = _RAND_603[15:0];
  _RAND_604 = {1{`RANDOM}};
  io_output_2_sr_15 = _RAND_604[15:0];
  _RAND_605 = {1{`RANDOM}};
  io_output_2_sr_16 = _RAND_605[15:0];
  _RAND_606 = {1{`RANDOM}};
  io_output_2_sr_17 = _RAND_606[15:0];
  _RAND_607 = {1{`RANDOM}};
  io_output_2_sr_18 = _RAND_607[15:0];
  _RAND_608 = {1{`RANDOM}};
  io_output_2_sr_19 = _RAND_608[15:0];
  _RAND_609 = {1{`RANDOM}};
  io_output_2_sr_20 = _RAND_609[15:0];
  _RAND_610 = {1{`RANDOM}};
  io_output_2_sr_21 = _RAND_610[15:0];
  _RAND_611 = {1{`RANDOM}};
  io_output_2_sr_22 = _RAND_611[15:0];
  _RAND_612 = {1{`RANDOM}};
  io_output_2_sr_23 = _RAND_612[15:0];
  _RAND_613 = {1{`RANDOM}};
  io_output_2_sr_24 = _RAND_613[15:0];
  _RAND_614 = {1{`RANDOM}};
  io_output_2_sr_25 = _RAND_614[15:0];
  _RAND_615 = {1{`RANDOM}};
  io_output_2_sr_26 = _RAND_615[15:0];
  _RAND_616 = {1{`RANDOM}};
  io_output_2_sr_27 = _RAND_616[15:0];
  _RAND_617 = {1{`RANDOM}};
  io_output_2_sr_28 = _RAND_617[15:0];
  _RAND_618 = {1{`RANDOM}};
  io_output_3_sr_0 = _RAND_618[15:0];
  _RAND_619 = {1{`RANDOM}};
  io_output_3_sr_1 = _RAND_619[15:0];
  _RAND_620 = {1{`RANDOM}};
  io_output_3_sr_2 = _RAND_620[15:0];
  _RAND_621 = {1{`RANDOM}};
  io_output_3_sr_3 = _RAND_621[15:0];
  _RAND_622 = {1{`RANDOM}};
  io_output_3_sr_4 = _RAND_622[15:0];
  _RAND_623 = {1{`RANDOM}};
  io_output_3_sr_5 = _RAND_623[15:0];
  _RAND_624 = {1{`RANDOM}};
  io_output_3_sr_6 = _RAND_624[15:0];
  _RAND_625 = {1{`RANDOM}};
  io_output_3_sr_7 = _RAND_625[15:0];
  _RAND_626 = {1{`RANDOM}};
  io_output_3_sr_8 = _RAND_626[15:0];
  _RAND_627 = {1{`RANDOM}};
  io_output_3_sr_9 = _RAND_627[15:0];
  _RAND_628 = {1{`RANDOM}};
  io_output_3_sr_10 = _RAND_628[15:0];
  _RAND_629 = {1{`RANDOM}};
  io_output_3_sr_11 = _RAND_629[15:0];
  _RAND_630 = {1{`RANDOM}};
  io_output_3_sr_12 = _RAND_630[15:0];
  _RAND_631 = {1{`RANDOM}};
  io_output_3_sr_13 = _RAND_631[15:0];
  _RAND_632 = {1{`RANDOM}};
  io_output_3_sr_14 = _RAND_632[15:0];
  _RAND_633 = {1{`RANDOM}};
  io_output_3_sr_15 = _RAND_633[15:0];
  _RAND_634 = {1{`RANDOM}};
  io_output_3_sr_16 = _RAND_634[15:0];
  _RAND_635 = {1{`RANDOM}};
  io_output_3_sr_17 = _RAND_635[15:0];
  _RAND_636 = {1{`RANDOM}};
  io_output_3_sr_18 = _RAND_636[15:0];
  _RAND_637 = {1{`RANDOM}};
  io_output_3_sr_19 = _RAND_637[15:0];
  _RAND_638 = {1{`RANDOM}};
  io_output_3_sr_20 = _RAND_638[15:0];
  _RAND_639 = {1{`RANDOM}};
  io_output_3_sr_21 = _RAND_639[15:0];
  _RAND_640 = {1{`RANDOM}};
  io_output_3_sr_22 = _RAND_640[15:0];
  _RAND_641 = {1{`RANDOM}};
  io_output_3_sr_23 = _RAND_641[15:0];
  _RAND_642 = {1{`RANDOM}};
  io_output_3_sr_24 = _RAND_642[15:0];
  _RAND_643 = {1{`RANDOM}};
  io_output_3_sr_25 = _RAND_643[15:0];
  _RAND_644 = {1{`RANDOM}};
  io_output_3_sr_26 = _RAND_644[15:0];
  _RAND_645 = {1{`RANDOM}};
  io_output_3_sr_27 = _RAND_645[15:0];
  _RAND_646 = {1{`RANDOM}};
  io_output_4_sr_0 = _RAND_646[15:0];
  _RAND_647 = {1{`RANDOM}};
  io_output_4_sr_1 = _RAND_647[15:0];
  _RAND_648 = {1{`RANDOM}};
  io_output_4_sr_2 = _RAND_648[15:0];
  _RAND_649 = {1{`RANDOM}};
  io_output_4_sr_3 = _RAND_649[15:0];
  _RAND_650 = {1{`RANDOM}};
  io_output_4_sr_4 = _RAND_650[15:0];
  _RAND_651 = {1{`RANDOM}};
  io_output_4_sr_5 = _RAND_651[15:0];
  _RAND_652 = {1{`RANDOM}};
  io_output_4_sr_6 = _RAND_652[15:0];
  _RAND_653 = {1{`RANDOM}};
  io_output_4_sr_7 = _RAND_653[15:0];
  _RAND_654 = {1{`RANDOM}};
  io_output_4_sr_8 = _RAND_654[15:0];
  _RAND_655 = {1{`RANDOM}};
  io_output_4_sr_9 = _RAND_655[15:0];
  _RAND_656 = {1{`RANDOM}};
  io_output_4_sr_10 = _RAND_656[15:0];
  _RAND_657 = {1{`RANDOM}};
  io_output_4_sr_11 = _RAND_657[15:0];
  _RAND_658 = {1{`RANDOM}};
  io_output_4_sr_12 = _RAND_658[15:0];
  _RAND_659 = {1{`RANDOM}};
  io_output_4_sr_13 = _RAND_659[15:0];
  _RAND_660 = {1{`RANDOM}};
  io_output_4_sr_14 = _RAND_660[15:0];
  _RAND_661 = {1{`RANDOM}};
  io_output_4_sr_15 = _RAND_661[15:0];
  _RAND_662 = {1{`RANDOM}};
  io_output_4_sr_16 = _RAND_662[15:0];
  _RAND_663 = {1{`RANDOM}};
  io_output_4_sr_17 = _RAND_663[15:0];
  _RAND_664 = {1{`RANDOM}};
  io_output_4_sr_18 = _RAND_664[15:0];
  _RAND_665 = {1{`RANDOM}};
  io_output_4_sr_19 = _RAND_665[15:0];
  _RAND_666 = {1{`RANDOM}};
  io_output_4_sr_20 = _RAND_666[15:0];
  _RAND_667 = {1{`RANDOM}};
  io_output_4_sr_21 = _RAND_667[15:0];
  _RAND_668 = {1{`RANDOM}};
  io_output_4_sr_22 = _RAND_668[15:0];
  _RAND_669 = {1{`RANDOM}};
  io_output_4_sr_23 = _RAND_669[15:0];
  _RAND_670 = {1{`RANDOM}};
  io_output_4_sr_24 = _RAND_670[15:0];
  _RAND_671 = {1{`RANDOM}};
  io_output_4_sr_25 = _RAND_671[15:0];
  _RAND_672 = {1{`RANDOM}};
  io_output_4_sr_26 = _RAND_672[15:0];
  _RAND_673 = {1{`RANDOM}};
  io_output_5_sr_0 = _RAND_673[15:0];
  _RAND_674 = {1{`RANDOM}};
  io_output_5_sr_1 = _RAND_674[15:0];
  _RAND_675 = {1{`RANDOM}};
  io_output_5_sr_2 = _RAND_675[15:0];
  _RAND_676 = {1{`RANDOM}};
  io_output_5_sr_3 = _RAND_676[15:0];
  _RAND_677 = {1{`RANDOM}};
  io_output_5_sr_4 = _RAND_677[15:0];
  _RAND_678 = {1{`RANDOM}};
  io_output_5_sr_5 = _RAND_678[15:0];
  _RAND_679 = {1{`RANDOM}};
  io_output_5_sr_6 = _RAND_679[15:0];
  _RAND_680 = {1{`RANDOM}};
  io_output_5_sr_7 = _RAND_680[15:0];
  _RAND_681 = {1{`RANDOM}};
  io_output_5_sr_8 = _RAND_681[15:0];
  _RAND_682 = {1{`RANDOM}};
  io_output_5_sr_9 = _RAND_682[15:0];
  _RAND_683 = {1{`RANDOM}};
  io_output_5_sr_10 = _RAND_683[15:0];
  _RAND_684 = {1{`RANDOM}};
  io_output_5_sr_11 = _RAND_684[15:0];
  _RAND_685 = {1{`RANDOM}};
  io_output_5_sr_12 = _RAND_685[15:0];
  _RAND_686 = {1{`RANDOM}};
  io_output_5_sr_13 = _RAND_686[15:0];
  _RAND_687 = {1{`RANDOM}};
  io_output_5_sr_14 = _RAND_687[15:0];
  _RAND_688 = {1{`RANDOM}};
  io_output_5_sr_15 = _RAND_688[15:0];
  _RAND_689 = {1{`RANDOM}};
  io_output_5_sr_16 = _RAND_689[15:0];
  _RAND_690 = {1{`RANDOM}};
  io_output_5_sr_17 = _RAND_690[15:0];
  _RAND_691 = {1{`RANDOM}};
  io_output_5_sr_18 = _RAND_691[15:0];
  _RAND_692 = {1{`RANDOM}};
  io_output_5_sr_19 = _RAND_692[15:0];
  _RAND_693 = {1{`RANDOM}};
  io_output_5_sr_20 = _RAND_693[15:0];
  _RAND_694 = {1{`RANDOM}};
  io_output_5_sr_21 = _RAND_694[15:0];
  _RAND_695 = {1{`RANDOM}};
  io_output_5_sr_22 = _RAND_695[15:0];
  _RAND_696 = {1{`RANDOM}};
  io_output_5_sr_23 = _RAND_696[15:0];
  _RAND_697 = {1{`RANDOM}};
  io_output_5_sr_24 = _RAND_697[15:0];
  _RAND_698 = {1{`RANDOM}};
  io_output_5_sr_25 = _RAND_698[15:0];
  _RAND_699 = {1{`RANDOM}};
  io_output_6_sr_0 = _RAND_699[15:0];
  _RAND_700 = {1{`RANDOM}};
  io_output_6_sr_1 = _RAND_700[15:0];
  _RAND_701 = {1{`RANDOM}};
  io_output_6_sr_2 = _RAND_701[15:0];
  _RAND_702 = {1{`RANDOM}};
  io_output_6_sr_3 = _RAND_702[15:0];
  _RAND_703 = {1{`RANDOM}};
  io_output_6_sr_4 = _RAND_703[15:0];
  _RAND_704 = {1{`RANDOM}};
  io_output_6_sr_5 = _RAND_704[15:0];
  _RAND_705 = {1{`RANDOM}};
  io_output_6_sr_6 = _RAND_705[15:0];
  _RAND_706 = {1{`RANDOM}};
  io_output_6_sr_7 = _RAND_706[15:0];
  _RAND_707 = {1{`RANDOM}};
  io_output_6_sr_8 = _RAND_707[15:0];
  _RAND_708 = {1{`RANDOM}};
  io_output_6_sr_9 = _RAND_708[15:0];
  _RAND_709 = {1{`RANDOM}};
  io_output_6_sr_10 = _RAND_709[15:0];
  _RAND_710 = {1{`RANDOM}};
  io_output_6_sr_11 = _RAND_710[15:0];
  _RAND_711 = {1{`RANDOM}};
  io_output_6_sr_12 = _RAND_711[15:0];
  _RAND_712 = {1{`RANDOM}};
  io_output_6_sr_13 = _RAND_712[15:0];
  _RAND_713 = {1{`RANDOM}};
  io_output_6_sr_14 = _RAND_713[15:0];
  _RAND_714 = {1{`RANDOM}};
  io_output_6_sr_15 = _RAND_714[15:0];
  _RAND_715 = {1{`RANDOM}};
  io_output_6_sr_16 = _RAND_715[15:0];
  _RAND_716 = {1{`RANDOM}};
  io_output_6_sr_17 = _RAND_716[15:0];
  _RAND_717 = {1{`RANDOM}};
  io_output_6_sr_18 = _RAND_717[15:0];
  _RAND_718 = {1{`RANDOM}};
  io_output_6_sr_19 = _RAND_718[15:0];
  _RAND_719 = {1{`RANDOM}};
  io_output_6_sr_20 = _RAND_719[15:0];
  _RAND_720 = {1{`RANDOM}};
  io_output_6_sr_21 = _RAND_720[15:0];
  _RAND_721 = {1{`RANDOM}};
  io_output_6_sr_22 = _RAND_721[15:0];
  _RAND_722 = {1{`RANDOM}};
  io_output_6_sr_23 = _RAND_722[15:0];
  _RAND_723 = {1{`RANDOM}};
  io_output_6_sr_24 = _RAND_723[15:0];
  _RAND_724 = {1{`RANDOM}};
  io_output_7_sr_0 = _RAND_724[15:0];
  _RAND_725 = {1{`RANDOM}};
  io_output_7_sr_1 = _RAND_725[15:0];
  _RAND_726 = {1{`RANDOM}};
  io_output_7_sr_2 = _RAND_726[15:0];
  _RAND_727 = {1{`RANDOM}};
  io_output_7_sr_3 = _RAND_727[15:0];
  _RAND_728 = {1{`RANDOM}};
  io_output_7_sr_4 = _RAND_728[15:0];
  _RAND_729 = {1{`RANDOM}};
  io_output_7_sr_5 = _RAND_729[15:0];
  _RAND_730 = {1{`RANDOM}};
  io_output_7_sr_6 = _RAND_730[15:0];
  _RAND_731 = {1{`RANDOM}};
  io_output_7_sr_7 = _RAND_731[15:0];
  _RAND_732 = {1{`RANDOM}};
  io_output_7_sr_8 = _RAND_732[15:0];
  _RAND_733 = {1{`RANDOM}};
  io_output_7_sr_9 = _RAND_733[15:0];
  _RAND_734 = {1{`RANDOM}};
  io_output_7_sr_10 = _RAND_734[15:0];
  _RAND_735 = {1{`RANDOM}};
  io_output_7_sr_11 = _RAND_735[15:0];
  _RAND_736 = {1{`RANDOM}};
  io_output_7_sr_12 = _RAND_736[15:0];
  _RAND_737 = {1{`RANDOM}};
  io_output_7_sr_13 = _RAND_737[15:0];
  _RAND_738 = {1{`RANDOM}};
  io_output_7_sr_14 = _RAND_738[15:0];
  _RAND_739 = {1{`RANDOM}};
  io_output_7_sr_15 = _RAND_739[15:0];
  _RAND_740 = {1{`RANDOM}};
  io_output_7_sr_16 = _RAND_740[15:0];
  _RAND_741 = {1{`RANDOM}};
  io_output_7_sr_17 = _RAND_741[15:0];
  _RAND_742 = {1{`RANDOM}};
  io_output_7_sr_18 = _RAND_742[15:0];
  _RAND_743 = {1{`RANDOM}};
  io_output_7_sr_19 = _RAND_743[15:0];
  _RAND_744 = {1{`RANDOM}};
  io_output_7_sr_20 = _RAND_744[15:0];
  _RAND_745 = {1{`RANDOM}};
  io_output_7_sr_21 = _RAND_745[15:0];
  _RAND_746 = {1{`RANDOM}};
  io_output_7_sr_22 = _RAND_746[15:0];
  _RAND_747 = {1{`RANDOM}};
  io_output_7_sr_23 = _RAND_747[15:0];
  _RAND_748 = {1{`RANDOM}};
  io_output_8_sr_0 = _RAND_748[15:0];
  _RAND_749 = {1{`RANDOM}};
  io_output_8_sr_1 = _RAND_749[15:0];
  _RAND_750 = {1{`RANDOM}};
  io_output_8_sr_2 = _RAND_750[15:0];
  _RAND_751 = {1{`RANDOM}};
  io_output_8_sr_3 = _RAND_751[15:0];
  _RAND_752 = {1{`RANDOM}};
  io_output_8_sr_4 = _RAND_752[15:0];
  _RAND_753 = {1{`RANDOM}};
  io_output_8_sr_5 = _RAND_753[15:0];
  _RAND_754 = {1{`RANDOM}};
  io_output_8_sr_6 = _RAND_754[15:0];
  _RAND_755 = {1{`RANDOM}};
  io_output_8_sr_7 = _RAND_755[15:0];
  _RAND_756 = {1{`RANDOM}};
  io_output_8_sr_8 = _RAND_756[15:0];
  _RAND_757 = {1{`RANDOM}};
  io_output_8_sr_9 = _RAND_757[15:0];
  _RAND_758 = {1{`RANDOM}};
  io_output_8_sr_10 = _RAND_758[15:0];
  _RAND_759 = {1{`RANDOM}};
  io_output_8_sr_11 = _RAND_759[15:0];
  _RAND_760 = {1{`RANDOM}};
  io_output_8_sr_12 = _RAND_760[15:0];
  _RAND_761 = {1{`RANDOM}};
  io_output_8_sr_13 = _RAND_761[15:0];
  _RAND_762 = {1{`RANDOM}};
  io_output_8_sr_14 = _RAND_762[15:0];
  _RAND_763 = {1{`RANDOM}};
  io_output_8_sr_15 = _RAND_763[15:0];
  _RAND_764 = {1{`RANDOM}};
  io_output_8_sr_16 = _RAND_764[15:0];
  _RAND_765 = {1{`RANDOM}};
  io_output_8_sr_17 = _RAND_765[15:0];
  _RAND_766 = {1{`RANDOM}};
  io_output_8_sr_18 = _RAND_766[15:0];
  _RAND_767 = {1{`RANDOM}};
  io_output_8_sr_19 = _RAND_767[15:0];
  _RAND_768 = {1{`RANDOM}};
  io_output_8_sr_20 = _RAND_768[15:0];
  _RAND_769 = {1{`RANDOM}};
  io_output_8_sr_21 = _RAND_769[15:0];
  _RAND_770 = {1{`RANDOM}};
  io_output_8_sr_22 = _RAND_770[15:0];
  _RAND_771 = {1{`RANDOM}};
  io_output_9_sr_0 = _RAND_771[15:0];
  _RAND_772 = {1{`RANDOM}};
  io_output_9_sr_1 = _RAND_772[15:0];
  _RAND_773 = {1{`RANDOM}};
  io_output_9_sr_2 = _RAND_773[15:0];
  _RAND_774 = {1{`RANDOM}};
  io_output_9_sr_3 = _RAND_774[15:0];
  _RAND_775 = {1{`RANDOM}};
  io_output_9_sr_4 = _RAND_775[15:0];
  _RAND_776 = {1{`RANDOM}};
  io_output_9_sr_5 = _RAND_776[15:0];
  _RAND_777 = {1{`RANDOM}};
  io_output_9_sr_6 = _RAND_777[15:0];
  _RAND_778 = {1{`RANDOM}};
  io_output_9_sr_7 = _RAND_778[15:0];
  _RAND_779 = {1{`RANDOM}};
  io_output_9_sr_8 = _RAND_779[15:0];
  _RAND_780 = {1{`RANDOM}};
  io_output_9_sr_9 = _RAND_780[15:0];
  _RAND_781 = {1{`RANDOM}};
  io_output_9_sr_10 = _RAND_781[15:0];
  _RAND_782 = {1{`RANDOM}};
  io_output_9_sr_11 = _RAND_782[15:0];
  _RAND_783 = {1{`RANDOM}};
  io_output_9_sr_12 = _RAND_783[15:0];
  _RAND_784 = {1{`RANDOM}};
  io_output_9_sr_13 = _RAND_784[15:0];
  _RAND_785 = {1{`RANDOM}};
  io_output_9_sr_14 = _RAND_785[15:0];
  _RAND_786 = {1{`RANDOM}};
  io_output_9_sr_15 = _RAND_786[15:0];
  _RAND_787 = {1{`RANDOM}};
  io_output_9_sr_16 = _RAND_787[15:0];
  _RAND_788 = {1{`RANDOM}};
  io_output_9_sr_17 = _RAND_788[15:0];
  _RAND_789 = {1{`RANDOM}};
  io_output_9_sr_18 = _RAND_789[15:0];
  _RAND_790 = {1{`RANDOM}};
  io_output_9_sr_19 = _RAND_790[15:0];
  _RAND_791 = {1{`RANDOM}};
  io_output_9_sr_20 = _RAND_791[15:0];
  _RAND_792 = {1{`RANDOM}};
  io_output_9_sr_21 = _RAND_792[15:0];
  _RAND_793 = {1{`RANDOM}};
  io_output_10_sr_0 = _RAND_793[15:0];
  _RAND_794 = {1{`RANDOM}};
  io_output_10_sr_1 = _RAND_794[15:0];
  _RAND_795 = {1{`RANDOM}};
  io_output_10_sr_2 = _RAND_795[15:0];
  _RAND_796 = {1{`RANDOM}};
  io_output_10_sr_3 = _RAND_796[15:0];
  _RAND_797 = {1{`RANDOM}};
  io_output_10_sr_4 = _RAND_797[15:0];
  _RAND_798 = {1{`RANDOM}};
  io_output_10_sr_5 = _RAND_798[15:0];
  _RAND_799 = {1{`RANDOM}};
  io_output_10_sr_6 = _RAND_799[15:0];
  _RAND_800 = {1{`RANDOM}};
  io_output_10_sr_7 = _RAND_800[15:0];
  _RAND_801 = {1{`RANDOM}};
  io_output_10_sr_8 = _RAND_801[15:0];
  _RAND_802 = {1{`RANDOM}};
  io_output_10_sr_9 = _RAND_802[15:0];
  _RAND_803 = {1{`RANDOM}};
  io_output_10_sr_10 = _RAND_803[15:0];
  _RAND_804 = {1{`RANDOM}};
  io_output_10_sr_11 = _RAND_804[15:0];
  _RAND_805 = {1{`RANDOM}};
  io_output_10_sr_12 = _RAND_805[15:0];
  _RAND_806 = {1{`RANDOM}};
  io_output_10_sr_13 = _RAND_806[15:0];
  _RAND_807 = {1{`RANDOM}};
  io_output_10_sr_14 = _RAND_807[15:0];
  _RAND_808 = {1{`RANDOM}};
  io_output_10_sr_15 = _RAND_808[15:0];
  _RAND_809 = {1{`RANDOM}};
  io_output_10_sr_16 = _RAND_809[15:0];
  _RAND_810 = {1{`RANDOM}};
  io_output_10_sr_17 = _RAND_810[15:0];
  _RAND_811 = {1{`RANDOM}};
  io_output_10_sr_18 = _RAND_811[15:0];
  _RAND_812 = {1{`RANDOM}};
  io_output_10_sr_19 = _RAND_812[15:0];
  _RAND_813 = {1{`RANDOM}};
  io_output_10_sr_20 = _RAND_813[15:0];
  _RAND_814 = {1{`RANDOM}};
  io_output_11_sr_0 = _RAND_814[15:0];
  _RAND_815 = {1{`RANDOM}};
  io_output_11_sr_1 = _RAND_815[15:0];
  _RAND_816 = {1{`RANDOM}};
  io_output_11_sr_2 = _RAND_816[15:0];
  _RAND_817 = {1{`RANDOM}};
  io_output_11_sr_3 = _RAND_817[15:0];
  _RAND_818 = {1{`RANDOM}};
  io_output_11_sr_4 = _RAND_818[15:0];
  _RAND_819 = {1{`RANDOM}};
  io_output_11_sr_5 = _RAND_819[15:0];
  _RAND_820 = {1{`RANDOM}};
  io_output_11_sr_6 = _RAND_820[15:0];
  _RAND_821 = {1{`RANDOM}};
  io_output_11_sr_7 = _RAND_821[15:0];
  _RAND_822 = {1{`RANDOM}};
  io_output_11_sr_8 = _RAND_822[15:0];
  _RAND_823 = {1{`RANDOM}};
  io_output_11_sr_9 = _RAND_823[15:0];
  _RAND_824 = {1{`RANDOM}};
  io_output_11_sr_10 = _RAND_824[15:0];
  _RAND_825 = {1{`RANDOM}};
  io_output_11_sr_11 = _RAND_825[15:0];
  _RAND_826 = {1{`RANDOM}};
  io_output_11_sr_12 = _RAND_826[15:0];
  _RAND_827 = {1{`RANDOM}};
  io_output_11_sr_13 = _RAND_827[15:0];
  _RAND_828 = {1{`RANDOM}};
  io_output_11_sr_14 = _RAND_828[15:0];
  _RAND_829 = {1{`RANDOM}};
  io_output_11_sr_15 = _RAND_829[15:0];
  _RAND_830 = {1{`RANDOM}};
  io_output_11_sr_16 = _RAND_830[15:0];
  _RAND_831 = {1{`RANDOM}};
  io_output_11_sr_17 = _RAND_831[15:0];
  _RAND_832 = {1{`RANDOM}};
  io_output_11_sr_18 = _RAND_832[15:0];
  _RAND_833 = {1{`RANDOM}};
  io_output_11_sr_19 = _RAND_833[15:0];
  _RAND_834 = {1{`RANDOM}};
  io_output_12_sr_0 = _RAND_834[15:0];
  _RAND_835 = {1{`RANDOM}};
  io_output_12_sr_1 = _RAND_835[15:0];
  _RAND_836 = {1{`RANDOM}};
  io_output_12_sr_2 = _RAND_836[15:0];
  _RAND_837 = {1{`RANDOM}};
  io_output_12_sr_3 = _RAND_837[15:0];
  _RAND_838 = {1{`RANDOM}};
  io_output_12_sr_4 = _RAND_838[15:0];
  _RAND_839 = {1{`RANDOM}};
  io_output_12_sr_5 = _RAND_839[15:0];
  _RAND_840 = {1{`RANDOM}};
  io_output_12_sr_6 = _RAND_840[15:0];
  _RAND_841 = {1{`RANDOM}};
  io_output_12_sr_7 = _RAND_841[15:0];
  _RAND_842 = {1{`RANDOM}};
  io_output_12_sr_8 = _RAND_842[15:0];
  _RAND_843 = {1{`RANDOM}};
  io_output_12_sr_9 = _RAND_843[15:0];
  _RAND_844 = {1{`RANDOM}};
  io_output_12_sr_10 = _RAND_844[15:0];
  _RAND_845 = {1{`RANDOM}};
  io_output_12_sr_11 = _RAND_845[15:0];
  _RAND_846 = {1{`RANDOM}};
  io_output_12_sr_12 = _RAND_846[15:0];
  _RAND_847 = {1{`RANDOM}};
  io_output_12_sr_13 = _RAND_847[15:0];
  _RAND_848 = {1{`RANDOM}};
  io_output_12_sr_14 = _RAND_848[15:0];
  _RAND_849 = {1{`RANDOM}};
  io_output_12_sr_15 = _RAND_849[15:0];
  _RAND_850 = {1{`RANDOM}};
  io_output_12_sr_16 = _RAND_850[15:0];
  _RAND_851 = {1{`RANDOM}};
  io_output_12_sr_17 = _RAND_851[15:0];
  _RAND_852 = {1{`RANDOM}};
  io_output_12_sr_18 = _RAND_852[15:0];
  _RAND_853 = {1{`RANDOM}};
  io_output_13_sr_0 = _RAND_853[15:0];
  _RAND_854 = {1{`RANDOM}};
  io_output_13_sr_1 = _RAND_854[15:0];
  _RAND_855 = {1{`RANDOM}};
  io_output_13_sr_2 = _RAND_855[15:0];
  _RAND_856 = {1{`RANDOM}};
  io_output_13_sr_3 = _RAND_856[15:0];
  _RAND_857 = {1{`RANDOM}};
  io_output_13_sr_4 = _RAND_857[15:0];
  _RAND_858 = {1{`RANDOM}};
  io_output_13_sr_5 = _RAND_858[15:0];
  _RAND_859 = {1{`RANDOM}};
  io_output_13_sr_6 = _RAND_859[15:0];
  _RAND_860 = {1{`RANDOM}};
  io_output_13_sr_7 = _RAND_860[15:0];
  _RAND_861 = {1{`RANDOM}};
  io_output_13_sr_8 = _RAND_861[15:0];
  _RAND_862 = {1{`RANDOM}};
  io_output_13_sr_9 = _RAND_862[15:0];
  _RAND_863 = {1{`RANDOM}};
  io_output_13_sr_10 = _RAND_863[15:0];
  _RAND_864 = {1{`RANDOM}};
  io_output_13_sr_11 = _RAND_864[15:0];
  _RAND_865 = {1{`RANDOM}};
  io_output_13_sr_12 = _RAND_865[15:0];
  _RAND_866 = {1{`RANDOM}};
  io_output_13_sr_13 = _RAND_866[15:0];
  _RAND_867 = {1{`RANDOM}};
  io_output_13_sr_14 = _RAND_867[15:0];
  _RAND_868 = {1{`RANDOM}};
  io_output_13_sr_15 = _RAND_868[15:0];
  _RAND_869 = {1{`RANDOM}};
  io_output_13_sr_16 = _RAND_869[15:0];
  _RAND_870 = {1{`RANDOM}};
  io_output_13_sr_17 = _RAND_870[15:0];
  _RAND_871 = {1{`RANDOM}};
  io_output_14_sr_0 = _RAND_871[15:0];
  _RAND_872 = {1{`RANDOM}};
  io_output_14_sr_1 = _RAND_872[15:0];
  _RAND_873 = {1{`RANDOM}};
  io_output_14_sr_2 = _RAND_873[15:0];
  _RAND_874 = {1{`RANDOM}};
  io_output_14_sr_3 = _RAND_874[15:0];
  _RAND_875 = {1{`RANDOM}};
  io_output_14_sr_4 = _RAND_875[15:0];
  _RAND_876 = {1{`RANDOM}};
  io_output_14_sr_5 = _RAND_876[15:0];
  _RAND_877 = {1{`RANDOM}};
  io_output_14_sr_6 = _RAND_877[15:0];
  _RAND_878 = {1{`RANDOM}};
  io_output_14_sr_7 = _RAND_878[15:0];
  _RAND_879 = {1{`RANDOM}};
  io_output_14_sr_8 = _RAND_879[15:0];
  _RAND_880 = {1{`RANDOM}};
  io_output_14_sr_9 = _RAND_880[15:0];
  _RAND_881 = {1{`RANDOM}};
  io_output_14_sr_10 = _RAND_881[15:0];
  _RAND_882 = {1{`RANDOM}};
  io_output_14_sr_11 = _RAND_882[15:0];
  _RAND_883 = {1{`RANDOM}};
  io_output_14_sr_12 = _RAND_883[15:0];
  _RAND_884 = {1{`RANDOM}};
  io_output_14_sr_13 = _RAND_884[15:0];
  _RAND_885 = {1{`RANDOM}};
  io_output_14_sr_14 = _RAND_885[15:0];
  _RAND_886 = {1{`RANDOM}};
  io_output_14_sr_15 = _RAND_886[15:0];
  _RAND_887 = {1{`RANDOM}};
  io_output_14_sr_16 = _RAND_887[15:0];
  _RAND_888 = {1{`RANDOM}};
  io_output_15_sr_0 = _RAND_888[15:0];
  _RAND_889 = {1{`RANDOM}};
  io_output_15_sr_1 = _RAND_889[15:0];
  _RAND_890 = {1{`RANDOM}};
  io_output_15_sr_2 = _RAND_890[15:0];
  _RAND_891 = {1{`RANDOM}};
  io_output_15_sr_3 = _RAND_891[15:0];
  _RAND_892 = {1{`RANDOM}};
  io_output_15_sr_4 = _RAND_892[15:0];
  _RAND_893 = {1{`RANDOM}};
  io_output_15_sr_5 = _RAND_893[15:0];
  _RAND_894 = {1{`RANDOM}};
  io_output_15_sr_6 = _RAND_894[15:0];
  _RAND_895 = {1{`RANDOM}};
  io_output_15_sr_7 = _RAND_895[15:0];
  _RAND_896 = {1{`RANDOM}};
  io_output_15_sr_8 = _RAND_896[15:0];
  _RAND_897 = {1{`RANDOM}};
  io_output_15_sr_9 = _RAND_897[15:0];
  _RAND_898 = {1{`RANDOM}};
  io_output_15_sr_10 = _RAND_898[15:0];
  _RAND_899 = {1{`RANDOM}};
  io_output_15_sr_11 = _RAND_899[15:0];
  _RAND_900 = {1{`RANDOM}};
  io_output_15_sr_12 = _RAND_900[15:0];
  _RAND_901 = {1{`RANDOM}};
  io_output_15_sr_13 = _RAND_901[15:0];
  _RAND_902 = {1{`RANDOM}};
  io_output_15_sr_14 = _RAND_902[15:0];
  _RAND_903 = {1{`RANDOM}};
  io_output_15_sr_15 = _RAND_903[15:0];
  _RAND_904 = {1{`RANDOM}};
  io_output_16_sr_0 = _RAND_904[15:0];
  _RAND_905 = {1{`RANDOM}};
  io_output_16_sr_1 = _RAND_905[15:0];
  _RAND_906 = {1{`RANDOM}};
  io_output_16_sr_2 = _RAND_906[15:0];
  _RAND_907 = {1{`RANDOM}};
  io_output_16_sr_3 = _RAND_907[15:0];
  _RAND_908 = {1{`RANDOM}};
  io_output_16_sr_4 = _RAND_908[15:0];
  _RAND_909 = {1{`RANDOM}};
  io_output_16_sr_5 = _RAND_909[15:0];
  _RAND_910 = {1{`RANDOM}};
  io_output_16_sr_6 = _RAND_910[15:0];
  _RAND_911 = {1{`RANDOM}};
  io_output_16_sr_7 = _RAND_911[15:0];
  _RAND_912 = {1{`RANDOM}};
  io_output_16_sr_8 = _RAND_912[15:0];
  _RAND_913 = {1{`RANDOM}};
  io_output_16_sr_9 = _RAND_913[15:0];
  _RAND_914 = {1{`RANDOM}};
  io_output_16_sr_10 = _RAND_914[15:0];
  _RAND_915 = {1{`RANDOM}};
  io_output_16_sr_11 = _RAND_915[15:0];
  _RAND_916 = {1{`RANDOM}};
  io_output_16_sr_12 = _RAND_916[15:0];
  _RAND_917 = {1{`RANDOM}};
  io_output_16_sr_13 = _RAND_917[15:0];
  _RAND_918 = {1{`RANDOM}};
  io_output_16_sr_14 = _RAND_918[15:0];
  _RAND_919 = {1{`RANDOM}};
  io_output_17_sr_0 = _RAND_919[15:0];
  _RAND_920 = {1{`RANDOM}};
  io_output_17_sr_1 = _RAND_920[15:0];
  _RAND_921 = {1{`RANDOM}};
  io_output_17_sr_2 = _RAND_921[15:0];
  _RAND_922 = {1{`RANDOM}};
  io_output_17_sr_3 = _RAND_922[15:0];
  _RAND_923 = {1{`RANDOM}};
  io_output_17_sr_4 = _RAND_923[15:0];
  _RAND_924 = {1{`RANDOM}};
  io_output_17_sr_5 = _RAND_924[15:0];
  _RAND_925 = {1{`RANDOM}};
  io_output_17_sr_6 = _RAND_925[15:0];
  _RAND_926 = {1{`RANDOM}};
  io_output_17_sr_7 = _RAND_926[15:0];
  _RAND_927 = {1{`RANDOM}};
  io_output_17_sr_8 = _RAND_927[15:0];
  _RAND_928 = {1{`RANDOM}};
  io_output_17_sr_9 = _RAND_928[15:0];
  _RAND_929 = {1{`RANDOM}};
  io_output_17_sr_10 = _RAND_929[15:0];
  _RAND_930 = {1{`RANDOM}};
  io_output_17_sr_11 = _RAND_930[15:0];
  _RAND_931 = {1{`RANDOM}};
  io_output_17_sr_12 = _RAND_931[15:0];
  _RAND_932 = {1{`RANDOM}};
  io_output_17_sr_13 = _RAND_932[15:0];
  _RAND_933 = {1{`RANDOM}};
  io_output_18_sr_0 = _RAND_933[15:0];
  _RAND_934 = {1{`RANDOM}};
  io_output_18_sr_1 = _RAND_934[15:0];
  _RAND_935 = {1{`RANDOM}};
  io_output_18_sr_2 = _RAND_935[15:0];
  _RAND_936 = {1{`RANDOM}};
  io_output_18_sr_3 = _RAND_936[15:0];
  _RAND_937 = {1{`RANDOM}};
  io_output_18_sr_4 = _RAND_937[15:0];
  _RAND_938 = {1{`RANDOM}};
  io_output_18_sr_5 = _RAND_938[15:0];
  _RAND_939 = {1{`RANDOM}};
  io_output_18_sr_6 = _RAND_939[15:0];
  _RAND_940 = {1{`RANDOM}};
  io_output_18_sr_7 = _RAND_940[15:0];
  _RAND_941 = {1{`RANDOM}};
  io_output_18_sr_8 = _RAND_941[15:0];
  _RAND_942 = {1{`RANDOM}};
  io_output_18_sr_9 = _RAND_942[15:0];
  _RAND_943 = {1{`RANDOM}};
  io_output_18_sr_10 = _RAND_943[15:0];
  _RAND_944 = {1{`RANDOM}};
  io_output_18_sr_11 = _RAND_944[15:0];
  _RAND_945 = {1{`RANDOM}};
  io_output_18_sr_12 = _RAND_945[15:0];
  _RAND_946 = {1{`RANDOM}};
  io_output_19_sr_0 = _RAND_946[15:0];
  _RAND_947 = {1{`RANDOM}};
  io_output_19_sr_1 = _RAND_947[15:0];
  _RAND_948 = {1{`RANDOM}};
  io_output_19_sr_2 = _RAND_948[15:0];
  _RAND_949 = {1{`RANDOM}};
  io_output_19_sr_3 = _RAND_949[15:0];
  _RAND_950 = {1{`RANDOM}};
  io_output_19_sr_4 = _RAND_950[15:0];
  _RAND_951 = {1{`RANDOM}};
  io_output_19_sr_5 = _RAND_951[15:0];
  _RAND_952 = {1{`RANDOM}};
  io_output_19_sr_6 = _RAND_952[15:0];
  _RAND_953 = {1{`RANDOM}};
  io_output_19_sr_7 = _RAND_953[15:0];
  _RAND_954 = {1{`RANDOM}};
  io_output_19_sr_8 = _RAND_954[15:0];
  _RAND_955 = {1{`RANDOM}};
  io_output_19_sr_9 = _RAND_955[15:0];
  _RAND_956 = {1{`RANDOM}};
  io_output_19_sr_10 = _RAND_956[15:0];
  _RAND_957 = {1{`RANDOM}};
  io_output_19_sr_11 = _RAND_957[15:0];
  _RAND_958 = {1{`RANDOM}};
  io_output_20_sr_0 = _RAND_958[15:0];
  _RAND_959 = {1{`RANDOM}};
  io_output_20_sr_1 = _RAND_959[15:0];
  _RAND_960 = {1{`RANDOM}};
  io_output_20_sr_2 = _RAND_960[15:0];
  _RAND_961 = {1{`RANDOM}};
  io_output_20_sr_3 = _RAND_961[15:0];
  _RAND_962 = {1{`RANDOM}};
  io_output_20_sr_4 = _RAND_962[15:0];
  _RAND_963 = {1{`RANDOM}};
  io_output_20_sr_5 = _RAND_963[15:0];
  _RAND_964 = {1{`RANDOM}};
  io_output_20_sr_6 = _RAND_964[15:0];
  _RAND_965 = {1{`RANDOM}};
  io_output_20_sr_7 = _RAND_965[15:0];
  _RAND_966 = {1{`RANDOM}};
  io_output_20_sr_8 = _RAND_966[15:0];
  _RAND_967 = {1{`RANDOM}};
  io_output_20_sr_9 = _RAND_967[15:0];
  _RAND_968 = {1{`RANDOM}};
  io_output_20_sr_10 = _RAND_968[15:0];
  _RAND_969 = {1{`RANDOM}};
  io_output_21_sr_0 = _RAND_969[15:0];
  _RAND_970 = {1{`RANDOM}};
  io_output_21_sr_1 = _RAND_970[15:0];
  _RAND_971 = {1{`RANDOM}};
  io_output_21_sr_2 = _RAND_971[15:0];
  _RAND_972 = {1{`RANDOM}};
  io_output_21_sr_3 = _RAND_972[15:0];
  _RAND_973 = {1{`RANDOM}};
  io_output_21_sr_4 = _RAND_973[15:0];
  _RAND_974 = {1{`RANDOM}};
  io_output_21_sr_5 = _RAND_974[15:0];
  _RAND_975 = {1{`RANDOM}};
  io_output_21_sr_6 = _RAND_975[15:0];
  _RAND_976 = {1{`RANDOM}};
  io_output_21_sr_7 = _RAND_976[15:0];
  _RAND_977 = {1{`RANDOM}};
  io_output_21_sr_8 = _RAND_977[15:0];
  _RAND_978 = {1{`RANDOM}};
  io_output_21_sr_9 = _RAND_978[15:0];
  _RAND_979 = {1{`RANDOM}};
  io_output_22_sr_0 = _RAND_979[15:0];
  _RAND_980 = {1{`RANDOM}};
  io_output_22_sr_1 = _RAND_980[15:0];
  _RAND_981 = {1{`RANDOM}};
  io_output_22_sr_2 = _RAND_981[15:0];
  _RAND_982 = {1{`RANDOM}};
  io_output_22_sr_3 = _RAND_982[15:0];
  _RAND_983 = {1{`RANDOM}};
  io_output_22_sr_4 = _RAND_983[15:0];
  _RAND_984 = {1{`RANDOM}};
  io_output_22_sr_5 = _RAND_984[15:0];
  _RAND_985 = {1{`RANDOM}};
  io_output_22_sr_6 = _RAND_985[15:0];
  _RAND_986 = {1{`RANDOM}};
  io_output_22_sr_7 = _RAND_986[15:0];
  _RAND_987 = {1{`RANDOM}};
  io_output_22_sr_8 = _RAND_987[15:0];
  _RAND_988 = {1{`RANDOM}};
  io_output_23_sr_0 = _RAND_988[15:0];
  _RAND_989 = {1{`RANDOM}};
  io_output_23_sr_1 = _RAND_989[15:0];
  _RAND_990 = {1{`RANDOM}};
  io_output_23_sr_2 = _RAND_990[15:0];
  _RAND_991 = {1{`RANDOM}};
  io_output_23_sr_3 = _RAND_991[15:0];
  _RAND_992 = {1{`RANDOM}};
  io_output_23_sr_4 = _RAND_992[15:0];
  _RAND_993 = {1{`RANDOM}};
  io_output_23_sr_5 = _RAND_993[15:0];
  _RAND_994 = {1{`RANDOM}};
  io_output_23_sr_6 = _RAND_994[15:0];
  _RAND_995 = {1{`RANDOM}};
  io_output_23_sr_7 = _RAND_995[15:0];
  _RAND_996 = {1{`RANDOM}};
  io_output_24_sr_0 = _RAND_996[15:0];
  _RAND_997 = {1{`RANDOM}};
  io_output_24_sr_1 = _RAND_997[15:0];
  _RAND_998 = {1{`RANDOM}};
  io_output_24_sr_2 = _RAND_998[15:0];
  _RAND_999 = {1{`RANDOM}};
  io_output_24_sr_3 = _RAND_999[15:0];
  _RAND_1000 = {1{`RANDOM}};
  io_output_24_sr_4 = _RAND_1000[15:0];
  _RAND_1001 = {1{`RANDOM}};
  io_output_24_sr_5 = _RAND_1001[15:0];
  _RAND_1002 = {1{`RANDOM}};
  io_output_24_sr_6 = _RAND_1002[15:0];
  _RAND_1003 = {1{`RANDOM}};
  io_output_25_sr_0 = _RAND_1003[15:0];
  _RAND_1004 = {1{`RANDOM}};
  io_output_25_sr_1 = _RAND_1004[15:0];
  _RAND_1005 = {1{`RANDOM}};
  io_output_25_sr_2 = _RAND_1005[15:0];
  _RAND_1006 = {1{`RANDOM}};
  io_output_25_sr_3 = _RAND_1006[15:0];
  _RAND_1007 = {1{`RANDOM}};
  io_output_25_sr_4 = _RAND_1007[15:0];
  _RAND_1008 = {1{`RANDOM}};
  io_output_25_sr_5 = _RAND_1008[15:0];
  _RAND_1009 = {1{`RANDOM}};
  io_output_26_sr_0 = _RAND_1009[15:0];
  _RAND_1010 = {1{`RANDOM}};
  io_output_26_sr_1 = _RAND_1010[15:0];
  _RAND_1011 = {1{`RANDOM}};
  io_output_26_sr_2 = _RAND_1011[15:0];
  _RAND_1012 = {1{`RANDOM}};
  io_output_26_sr_3 = _RAND_1012[15:0];
  _RAND_1013 = {1{`RANDOM}};
  io_output_26_sr_4 = _RAND_1013[15:0];
  _RAND_1014 = {1{`RANDOM}};
  io_output_27_sr_0 = _RAND_1014[15:0];
  _RAND_1015 = {1{`RANDOM}};
  io_output_27_sr_1 = _RAND_1015[15:0];
  _RAND_1016 = {1{`RANDOM}};
  io_output_27_sr_2 = _RAND_1016[15:0];
  _RAND_1017 = {1{`RANDOM}};
  io_output_27_sr_3 = _RAND_1017[15:0];
  _RAND_1018 = {1{`RANDOM}};
  io_output_28_sr_0 = _RAND_1018[15:0];
  _RAND_1019 = {1{`RANDOM}};
  io_output_28_sr_1 = _RAND_1019[15:0];
  _RAND_1020 = {1{`RANDOM}};
  io_output_28_sr_2 = _RAND_1020[15:0];
  _RAND_1021 = {1{`RANDOM}};
  io_output_29_sr_0 = _RAND_1021[15:0];
  _RAND_1022 = {1{`RANDOM}};
  io_output_29_sr_1 = _RAND_1022[15:0];
  _RAND_1023 = {1{`RANDOM}};
  io_output_30_sr_0 = _RAND_1023[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_0,
  input  [15:0] io_enq_bits_1,
  input  [15:0] io_enq_bits_2,
  input  [15:0] io_enq_bits_3,
  input  [15:0] io_enq_bits_4,
  input  [15:0] io_enq_bits_5,
  input  [15:0] io_enq_bits_6,
  input  [15:0] io_enq_bits_7,
  input  [15:0] io_enq_bits_8,
  input  [15:0] io_enq_bits_9,
  input  [15:0] io_enq_bits_10,
  input  [15:0] io_enq_bits_11,
  input  [15:0] io_enq_bits_12,
  input  [15:0] io_enq_bits_13,
  input  [15:0] io_enq_bits_14,
  input  [15:0] io_enq_bits_15,
  input  [15:0] io_enq_bits_16,
  input  [15:0] io_enq_bits_17,
  input  [15:0] io_enq_bits_18,
  input  [15:0] io_enq_bits_19,
  input  [15:0] io_enq_bits_20,
  input  [15:0] io_enq_bits_21,
  input  [15:0] io_enq_bits_22,
  input  [15:0] io_enq_bits_23,
  input  [15:0] io_enq_bits_24,
  input  [15:0] io_enq_bits_25,
  input  [15:0] io_enq_bits_26,
  input  [15:0] io_enq_bits_27,
  input  [15:0] io_enq_bits_28,
  input  [15:0] io_enq_bits_29,
  input  [15:0] io_enq_bits_30,
  input  [15:0] io_enq_bits_31,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_0,
  output [15:0] io_deq_bits_1,
  output [15:0] io_deq_bits_2,
  output [15:0] io_deq_bits_3,
  output [15:0] io_deq_bits_4,
  output [15:0] io_deq_bits_5,
  output [15:0] io_deq_bits_6,
  output [15:0] io_deq_bits_7,
  output [15:0] io_deq_bits_8,
  output [15:0] io_deq_bits_9,
  output [15:0] io_deq_bits_10,
  output [15:0] io_deq_bits_11,
  output [15:0] io_deq_bits_12,
  output [15:0] io_deq_bits_13,
  output [15:0] io_deq_bits_14,
  output [15:0] io_deq_bits_15,
  output [15:0] io_deq_bits_16,
  output [15:0] io_deq_bits_17,
  output [15:0] io_deq_bits_18,
  output [15:0] io_deq_bits_19,
  output [15:0] io_deq_bits_20,
  output [15:0] io_deq_bits_21,
  output [15:0] io_deq_bits_22,
  output [15:0] io_deq_bits_23,
  output [15:0] io_deq_bits_24,
  output [15:0] io_deq_bits_25,
  output [15:0] io_deq_bits_26,
  output [15:0] io_deq_bits_27,
  output [15:0] io_deq_bits_28,
  output [15:0] io_deq_bits_29,
  output [15:0] io_deq_bits_30,
  output [15:0] io_deq_bits_31
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_62;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ram_0 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_1 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_2 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_3 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_4 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_5 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_6 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_7 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_8 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_8_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_8_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_8_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_8_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_8_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_8_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_8_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_9 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_9_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_9_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_9_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_9_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_9_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_9_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_9_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_10 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_10_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_10_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_10_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_10_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_10_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_10_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_10_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_11 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_11_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_11_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_11_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_11_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_11_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_11_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_11_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_12 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_12_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_12_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_12_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_12_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_12_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_12_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_12_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_13 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_13_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_13_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_13_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_13_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_13_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_13_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_13_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_14 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_14_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_14_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_14_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_14_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_14_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_14_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_14_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_15 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_15_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_15_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_15_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_15_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_15_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_15_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_15_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_16 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_16_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_16_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_16_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_16_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_16_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_16_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_16_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_17 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_17_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_17_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_17_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_17_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_17_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_17_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_17_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_18 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_18_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_18_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_18_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_18_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_18_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_18_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_18_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_19 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_19_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_19_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_19_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_19_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_19_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_19_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_19_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_20 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_20_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_20_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_20_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_20_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_20_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_20_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_20_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_21 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_21_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_21_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_21_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_21_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_21_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_21_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_21_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_22 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_22_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_22_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_22_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_22_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_22_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_22_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_22_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_23 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_23_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_23_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_23_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_23_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_23_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_23_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_23_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_24 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_24_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_24_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_24_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_24_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_24_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_24_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_24_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_25 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_25_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_25_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_25_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_25_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_25_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_25_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_25_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_26 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_26_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_26_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_26_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_26_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_26_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_26_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_26_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_27 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_27_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_27_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_27_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_27_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_27_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_27_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_27_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_28 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_28_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_28_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_28_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_28_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_28_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_28_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_28_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_29 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_29_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_29_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_29_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_29_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_29_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_29_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_29_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_30 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_30_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_30_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_30_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_30_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_30_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_30_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_30_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_31 [0:62]; // @[Decoupled.scala 259:95]
  wire  ram_31_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_31_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_31_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_31_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_31_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_31_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_31_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [5:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  wrap = enq_ptr_value == 6'h3e; // @[Counter.scala 74:24]
  wire [5:0] _value_T_1 = enq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire  _GEN_45 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_45 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  wrap_1 = deq_ptr_value == 6'h3e; // @[Counter.scala 74:24]
  wire [5:0] _value_T_3 = deq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_0_io_deq_bits_MPORT_data = ram_0[ram_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_0_io_deq_bits_MPORT_data = ram_0_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_1[15:0] :
    ram_0[ram_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_0_MPORT_data = io_enq_bits_0;
  assign ram_0_MPORT_addr = enq_ptr_value;
  assign ram_0_MPORT_mask = 1'h1;
  assign ram_0_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_1_io_deq_bits_MPORT_data = ram_1[ram_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_1_io_deq_bits_MPORT_data = ram_1_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_3[15:0] :
    ram_1[ram_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_1_MPORT_data = io_enq_bits_1;
  assign ram_1_MPORT_addr = enq_ptr_value;
  assign ram_1_MPORT_mask = 1'h1;
  assign ram_1_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_2_io_deq_bits_MPORT_data = ram_2[ram_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_2_io_deq_bits_MPORT_data = ram_2_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_5[15:0] :
    ram_2[ram_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_2_MPORT_data = io_enq_bits_2;
  assign ram_2_MPORT_addr = enq_ptr_value;
  assign ram_2_MPORT_mask = 1'h1;
  assign ram_2_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_3_io_deq_bits_MPORT_data = ram_3[ram_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_3_io_deq_bits_MPORT_data = ram_3_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_7[15:0] :
    ram_3[ram_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_3_MPORT_data = io_enq_bits_3;
  assign ram_3_MPORT_addr = enq_ptr_value;
  assign ram_3_MPORT_mask = 1'h1;
  assign ram_3_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_4_io_deq_bits_MPORT_data = ram_4[ram_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_4_io_deq_bits_MPORT_data = ram_4_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_9[15:0] :
    ram_4[ram_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_4_MPORT_data = io_enq_bits_4;
  assign ram_4_MPORT_addr = enq_ptr_value;
  assign ram_4_MPORT_mask = 1'h1;
  assign ram_4_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_5_io_deq_bits_MPORT_data = ram_5[ram_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_5_io_deq_bits_MPORT_data = ram_5_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_11[15:0] :
    ram_5[ram_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_5_MPORT_data = io_enq_bits_5;
  assign ram_5_MPORT_addr = enq_ptr_value;
  assign ram_5_MPORT_mask = 1'h1;
  assign ram_5_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_6_io_deq_bits_MPORT_data = ram_6[ram_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_6_io_deq_bits_MPORT_data = ram_6_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_13[15:0] :
    ram_6[ram_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_6_MPORT_data = io_enq_bits_6;
  assign ram_6_MPORT_addr = enq_ptr_value;
  assign ram_6_MPORT_mask = 1'h1;
  assign ram_6_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_7_io_deq_bits_MPORT_data = ram_7[ram_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_7_io_deq_bits_MPORT_data = ram_7_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_15[15:0] :
    ram_7[ram_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_7_MPORT_data = io_enq_bits_7;
  assign ram_7_MPORT_addr = enq_ptr_value;
  assign ram_7_MPORT_mask = 1'h1;
  assign ram_7_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_8_io_deq_bits_MPORT_en = 1'h1;
  assign ram_8_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_8_io_deq_bits_MPORT_data = ram_8[ram_8_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_8_io_deq_bits_MPORT_data = ram_8_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_17[15:0] :
    ram_8[ram_8_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_8_MPORT_data = io_enq_bits_8;
  assign ram_8_MPORT_addr = enq_ptr_value;
  assign ram_8_MPORT_mask = 1'h1;
  assign ram_8_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_9_io_deq_bits_MPORT_en = 1'h1;
  assign ram_9_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_9_io_deq_bits_MPORT_data = ram_9[ram_9_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_9_io_deq_bits_MPORT_data = ram_9_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_19[15:0] :
    ram_9[ram_9_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_9_MPORT_data = io_enq_bits_9;
  assign ram_9_MPORT_addr = enq_ptr_value;
  assign ram_9_MPORT_mask = 1'h1;
  assign ram_9_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_10_io_deq_bits_MPORT_en = 1'h1;
  assign ram_10_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_10_io_deq_bits_MPORT_data = ram_10[ram_10_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_10_io_deq_bits_MPORT_data = ram_10_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_21[15:0] :
    ram_10[ram_10_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_10_MPORT_data = io_enq_bits_10;
  assign ram_10_MPORT_addr = enq_ptr_value;
  assign ram_10_MPORT_mask = 1'h1;
  assign ram_10_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_11_io_deq_bits_MPORT_en = 1'h1;
  assign ram_11_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_11_io_deq_bits_MPORT_data = ram_11[ram_11_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_11_io_deq_bits_MPORT_data = ram_11_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_23[15:0] :
    ram_11[ram_11_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_11_MPORT_data = io_enq_bits_11;
  assign ram_11_MPORT_addr = enq_ptr_value;
  assign ram_11_MPORT_mask = 1'h1;
  assign ram_11_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_12_io_deq_bits_MPORT_en = 1'h1;
  assign ram_12_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_12_io_deq_bits_MPORT_data = ram_12[ram_12_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_12_io_deq_bits_MPORT_data = ram_12_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_25[15:0] :
    ram_12[ram_12_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_12_MPORT_data = io_enq_bits_12;
  assign ram_12_MPORT_addr = enq_ptr_value;
  assign ram_12_MPORT_mask = 1'h1;
  assign ram_12_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_13_io_deq_bits_MPORT_en = 1'h1;
  assign ram_13_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_13_io_deq_bits_MPORT_data = ram_13[ram_13_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_13_io_deq_bits_MPORT_data = ram_13_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_27[15:0] :
    ram_13[ram_13_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_13_MPORT_data = io_enq_bits_13;
  assign ram_13_MPORT_addr = enq_ptr_value;
  assign ram_13_MPORT_mask = 1'h1;
  assign ram_13_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_14_io_deq_bits_MPORT_en = 1'h1;
  assign ram_14_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_14_io_deq_bits_MPORT_data = ram_14[ram_14_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_14_io_deq_bits_MPORT_data = ram_14_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_29[15:0] :
    ram_14[ram_14_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_14_MPORT_data = io_enq_bits_14;
  assign ram_14_MPORT_addr = enq_ptr_value;
  assign ram_14_MPORT_mask = 1'h1;
  assign ram_14_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_15_io_deq_bits_MPORT_en = 1'h1;
  assign ram_15_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_15_io_deq_bits_MPORT_data = ram_15[ram_15_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_15_io_deq_bits_MPORT_data = ram_15_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_31[15:0] :
    ram_15[ram_15_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_15_MPORT_data = io_enq_bits_15;
  assign ram_15_MPORT_addr = enq_ptr_value;
  assign ram_15_MPORT_mask = 1'h1;
  assign ram_15_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_16_io_deq_bits_MPORT_en = 1'h1;
  assign ram_16_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_16_io_deq_bits_MPORT_data = ram_16[ram_16_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_16_io_deq_bits_MPORT_data = ram_16_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_33[15:0] :
    ram_16[ram_16_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_16_MPORT_data = io_enq_bits_16;
  assign ram_16_MPORT_addr = enq_ptr_value;
  assign ram_16_MPORT_mask = 1'h1;
  assign ram_16_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_17_io_deq_bits_MPORT_en = 1'h1;
  assign ram_17_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_17_io_deq_bits_MPORT_data = ram_17[ram_17_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_17_io_deq_bits_MPORT_data = ram_17_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_35[15:0] :
    ram_17[ram_17_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_17_MPORT_data = io_enq_bits_17;
  assign ram_17_MPORT_addr = enq_ptr_value;
  assign ram_17_MPORT_mask = 1'h1;
  assign ram_17_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_18_io_deq_bits_MPORT_en = 1'h1;
  assign ram_18_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_18_io_deq_bits_MPORT_data = ram_18[ram_18_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_18_io_deq_bits_MPORT_data = ram_18_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_37[15:0] :
    ram_18[ram_18_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_18_MPORT_data = io_enq_bits_18;
  assign ram_18_MPORT_addr = enq_ptr_value;
  assign ram_18_MPORT_mask = 1'h1;
  assign ram_18_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_19_io_deq_bits_MPORT_en = 1'h1;
  assign ram_19_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_19_io_deq_bits_MPORT_data = ram_19[ram_19_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_19_io_deq_bits_MPORT_data = ram_19_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_39[15:0] :
    ram_19[ram_19_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_19_MPORT_data = io_enq_bits_19;
  assign ram_19_MPORT_addr = enq_ptr_value;
  assign ram_19_MPORT_mask = 1'h1;
  assign ram_19_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_20_io_deq_bits_MPORT_en = 1'h1;
  assign ram_20_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_20_io_deq_bits_MPORT_data = ram_20[ram_20_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_20_io_deq_bits_MPORT_data = ram_20_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_41[15:0] :
    ram_20[ram_20_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_20_MPORT_data = io_enq_bits_20;
  assign ram_20_MPORT_addr = enq_ptr_value;
  assign ram_20_MPORT_mask = 1'h1;
  assign ram_20_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_21_io_deq_bits_MPORT_en = 1'h1;
  assign ram_21_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_21_io_deq_bits_MPORT_data = ram_21[ram_21_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_21_io_deq_bits_MPORT_data = ram_21_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_43[15:0] :
    ram_21[ram_21_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_21_MPORT_data = io_enq_bits_21;
  assign ram_21_MPORT_addr = enq_ptr_value;
  assign ram_21_MPORT_mask = 1'h1;
  assign ram_21_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_22_io_deq_bits_MPORT_en = 1'h1;
  assign ram_22_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_22_io_deq_bits_MPORT_data = ram_22[ram_22_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_22_io_deq_bits_MPORT_data = ram_22_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_45[15:0] :
    ram_22[ram_22_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_22_MPORT_data = io_enq_bits_22;
  assign ram_22_MPORT_addr = enq_ptr_value;
  assign ram_22_MPORT_mask = 1'h1;
  assign ram_22_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_23_io_deq_bits_MPORT_en = 1'h1;
  assign ram_23_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_23_io_deq_bits_MPORT_data = ram_23[ram_23_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_23_io_deq_bits_MPORT_data = ram_23_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_47[15:0] :
    ram_23[ram_23_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_23_MPORT_data = io_enq_bits_23;
  assign ram_23_MPORT_addr = enq_ptr_value;
  assign ram_23_MPORT_mask = 1'h1;
  assign ram_23_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_24_io_deq_bits_MPORT_en = 1'h1;
  assign ram_24_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_24_io_deq_bits_MPORT_data = ram_24[ram_24_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_24_io_deq_bits_MPORT_data = ram_24_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_49[15:0] :
    ram_24[ram_24_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_24_MPORT_data = io_enq_bits_24;
  assign ram_24_MPORT_addr = enq_ptr_value;
  assign ram_24_MPORT_mask = 1'h1;
  assign ram_24_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_25_io_deq_bits_MPORT_en = 1'h1;
  assign ram_25_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_25_io_deq_bits_MPORT_data = ram_25[ram_25_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_25_io_deq_bits_MPORT_data = ram_25_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_51[15:0] :
    ram_25[ram_25_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_25_MPORT_data = io_enq_bits_25;
  assign ram_25_MPORT_addr = enq_ptr_value;
  assign ram_25_MPORT_mask = 1'h1;
  assign ram_25_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_26_io_deq_bits_MPORT_en = 1'h1;
  assign ram_26_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_26_io_deq_bits_MPORT_data = ram_26[ram_26_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_26_io_deq_bits_MPORT_data = ram_26_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_53[15:0] :
    ram_26[ram_26_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_26_MPORT_data = io_enq_bits_26;
  assign ram_26_MPORT_addr = enq_ptr_value;
  assign ram_26_MPORT_mask = 1'h1;
  assign ram_26_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_27_io_deq_bits_MPORT_en = 1'h1;
  assign ram_27_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_27_io_deq_bits_MPORT_data = ram_27[ram_27_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_27_io_deq_bits_MPORT_data = ram_27_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_55[15:0] :
    ram_27[ram_27_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_27_MPORT_data = io_enq_bits_27;
  assign ram_27_MPORT_addr = enq_ptr_value;
  assign ram_27_MPORT_mask = 1'h1;
  assign ram_27_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_28_io_deq_bits_MPORT_en = 1'h1;
  assign ram_28_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_28_io_deq_bits_MPORT_data = ram_28[ram_28_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_28_io_deq_bits_MPORT_data = ram_28_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_57[15:0] :
    ram_28[ram_28_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_28_MPORT_data = io_enq_bits_28;
  assign ram_28_MPORT_addr = enq_ptr_value;
  assign ram_28_MPORT_mask = 1'h1;
  assign ram_28_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_29_io_deq_bits_MPORT_en = 1'h1;
  assign ram_29_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_29_io_deq_bits_MPORT_data = ram_29[ram_29_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_29_io_deq_bits_MPORT_data = ram_29_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_59[15:0] :
    ram_29[ram_29_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_29_MPORT_data = io_enq_bits_29;
  assign ram_29_MPORT_addr = enq_ptr_value;
  assign ram_29_MPORT_mask = 1'h1;
  assign ram_29_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_30_io_deq_bits_MPORT_en = 1'h1;
  assign ram_30_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_30_io_deq_bits_MPORT_data = ram_30[ram_30_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_30_io_deq_bits_MPORT_data = ram_30_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_61[15:0] :
    ram_30[ram_30_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_30_MPORT_data = io_enq_bits_30;
  assign ram_30_MPORT_addr = enq_ptr_value;
  assign ram_30_MPORT_mask = 1'h1;
  assign ram_30_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_31_io_deq_bits_MPORT_en = 1'h1;
  assign ram_31_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_31_io_deq_bits_MPORT_data = ram_31[ram_31_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_31_io_deq_bits_MPORT_data = ram_31_io_deq_bits_MPORT_addr >= 6'h3f ? _RAND_63[15:0] :
    ram_31[ram_31_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_31_MPORT_data = io_enq_bits_31;
  assign ram_31_MPORT_addr = enq_ptr_value;
  assign ram_31_MPORT_mask = 1'h1;
  assign ram_31_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_0 = empty ? $signed(io_enq_bits_0) : $signed(ram_0_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_1 = empty ? $signed(io_enq_bits_1) : $signed(ram_1_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_2 = empty ? $signed(io_enq_bits_2) : $signed(ram_2_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_3 = empty ? $signed(io_enq_bits_3) : $signed(ram_3_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_4 = empty ? $signed(io_enq_bits_4) : $signed(ram_4_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_5 = empty ? $signed(io_enq_bits_5) : $signed(ram_5_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_6 = empty ? $signed(io_enq_bits_6) : $signed(ram_6_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_7 = empty ? $signed(io_enq_bits_7) : $signed(ram_7_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_8 = empty ? $signed(io_enq_bits_8) : $signed(ram_8_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_9 = empty ? $signed(io_enq_bits_9) : $signed(ram_9_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_10 = empty ? $signed(io_enq_bits_10) : $signed(ram_10_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_11 = empty ? $signed(io_enq_bits_11) : $signed(ram_11_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_12 = empty ? $signed(io_enq_bits_12) : $signed(ram_12_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_13 = empty ? $signed(io_enq_bits_13) : $signed(ram_13_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_14 = empty ? $signed(io_enq_bits_14) : $signed(ram_14_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_15 = empty ? $signed(io_enq_bits_15) : $signed(ram_15_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_16 = empty ? $signed(io_enq_bits_16) : $signed(ram_16_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_17 = empty ? $signed(io_enq_bits_17) : $signed(ram_17_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_18 = empty ? $signed(io_enq_bits_18) : $signed(ram_18_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_19 = empty ? $signed(io_enq_bits_19) : $signed(ram_19_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_20 = empty ? $signed(io_enq_bits_20) : $signed(ram_20_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_21 = empty ? $signed(io_enq_bits_21) : $signed(ram_21_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_22 = empty ? $signed(io_enq_bits_22) : $signed(ram_22_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_23 = empty ? $signed(io_enq_bits_23) : $signed(ram_23_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_24 = empty ? $signed(io_enq_bits_24) : $signed(ram_24_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_25 = empty ? $signed(io_enq_bits_25) : $signed(ram_25_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_26 = empty ? $signed(io_enq_bits_26) : $signed(ram_26_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_27 = empty ? $signed(io_enq_bits_27) : $signed(ram_27_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_28 = empty ? $signed(io_enq_bits_28) : $signed(ram_28_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_29 = empty ? $signed(io_enq_bits_29) : $signed(ram_29_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_30 = empty ? $signed(io_enq_bits_30) : $signed(ram_30_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_31 = empty ? $signed(io_enq_bits_31) : $signed(ram_31_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_0_MPORT_en & ram_0_MPORT_mask) begin
      ram_0[ram_0_MPORT_addr] <= ram_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_1_MPORT_en & ram_1_MPORT_mask) begin
      ram_1[ram_1_MPORT_addr] <= ram_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_2_MPORT_en & ram_2_MPORT_mask) begin
      ram_2[ram_2_MPORT_addr] <= ram_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_3_MPORT_en & ram_3_MPORT_mask) begin
      ram_3[ram_3_MPORT_addr] <= ram_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_4_MPORT_en & ram_4_MPORT_mask) begin
      ram_4[ram_4_MPORT_addr] <= ram_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_5_MPORT_en & ram_5_MPORT_mask) begin
      ram_5[ram_5_MPORT_addr] <= ram_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_6_MPORT_en & ram_6_MPORT_mask) begin
      ram_6[ram_6_MPORT_addr] <= ram_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_7_MPORT_en & ram_7_MPORT_mask) begin
      ram_7[ram_7_MPORT_addr] <= ram_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_8_MPORT_en & ram_8_MPORT_mask) begin
      ram_8[ram_8_MPORT_addr] <= ram_8_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_9_MPORT_en & ram_9_MPORT_mask) begin
      ram_9[ram_9_MPORT_addr] <= ram_9_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_10_MPORT_en & ram_10_MPORT_mask) begin
      ram_10[ram_10_MPORT_addr] <= ram_10_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_11_MPORT_en & ram_11_MPORT_mask) begin
      ram_11[ram_11_MPORT_addr] <= ram_11_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_12_MPORT_en & ram_12_MPORT_mask) begin
      ram_12[ram_12_MPORT_addr] <= ram_12_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_13_MPORT_en & ram_13_MPORT_mask) begin
      ram_13[ram_13_MPORT_addr] <= ram_13_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_14_MPORT_en & ram_14_MPORT_mask) begin
      ram_14[ram_14_MPORT_addr] <= ram_14_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_15_MPORT_en & ram_15_MPORT_mask) begin
      ram_15[ram_15_MPORT_addr] <= ram_15_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_16_MPORT_en & ram_16_MPORT_mask) begin
      ram_16[ram_16_MPORT_addr] <= ram_16_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_17_MPORT_en & ram_17_MPORT_mask) begin
      ram_17[ram_17_MPORT_addr] <= ram_17_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_18_MPORT_en & ram_18_MPORT_mask) begin
      ram_18[ram_18_MPORT_addr] <= ram_18_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_19_MPORT_en & ram_19_MPORT_mask) begin
      ram_19[ram_19_MPORT_addr] <= ram_19_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_20_MPORT_en & ram_20_MPORT_mask) begin
      ram_20[ram_20_MPORT_addr] <= ram_20_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_21_MPORT_en & ram_21_MPORT_mask) begin
      ram_21[ram_21_MPORT_addr] <= ram_21_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_22_MPORT_en & ram_22_MPORT_mask) begin
      ram_22[ram_22_MPORT_addr] <= ram_22_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_23_MPORT_en & ram_23_MPORT_mask) begin
      ram_23[ram_23_MPORT_addr] <= ram_23_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_24_MPORT_en & ram_24_MPORT_mask) begin
      ram_24[ram_24_MPORT_addr] <= ram_24_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_25_MPORT_en & ram_25_MPORT_mask) begin
      ram_25[ram_25_MPORT_addr] <= ram_25_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_26_MPORT_en & ram_26_MPORT_mask) begin
      ram_26[ram_26_MPORT_addr] <= ram_26_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_27_MPORT_en & ram_27_MPORT_mask) begin
      ram_27[ram_27_MPORT_addr] <= ram_27_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_28_MPORT_en & ram_28_MPORT_mask) begin
      ram_28[ram_28_MPORT_addr] <= ram_28_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_29_MPORT_en & ram_29_MPORT_mask) begin
      ram_29[ram_29_MPORT_addr] <= ram_29_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_30_MPORT_en & ram_30_MPORT_mask) begin
      ram_30[ram_30_MPORT_addr] <= ram_30_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_31_MPORT_en & ram_31_MPORT_mask) begin
      ram_31[ram_31_MPORT_addr] <= ram_31_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      if (wrap) begin // @[Counter.scala 88:20]
        enq_ptr_value <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      if (wrap_1) begin // @[Counter.scala 88:20]
        deq_ptr_value <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
  _RAND_17 = {1{`RANDOM}};
  _RAND_19 = {1{`RANDOM}};
  _RAND_21 = {1{`RANDOM}};
  _RAND_23 = {1{`RANDOM}};
  _RAND_25 = {1{`RANDOM}};
  _RAND_27 = {1{`RANDOM}};
  _RAND_29 = {1{`RANDOM}};
  _RAND_31 = {1{`RANDOM}};
  _RAND_33 = {1{`RANDOM}};
  _RAND_35 = {1{`RANDOM}};
  _RAND_37 = {1{`RANDOM}};
  _RAND_39 = {1{`RANDOM}};
  _RAND_41 = {1{`RANDOM}};
  _RAND_43 = {1{`RANDOM}};
  _RAND_45 = {1{`RANDOM}};
  _RAND_47 = {1{`RANDOM}};
  _RAND_49 = {1{`RANDOM}};
  _RAND_51 = {1{`RANDOM}};
  _RAND_53 = {1{`RANDOM}};
  _RAND_55 = {1{`RANDOM}};
  _RAND_57 = {1{`RANDOM}};
  _RAND_59 = {1{`RANDOM}};
  _RAND_61 = {1{`RANDOM}};
  _RAND_63 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_0[initvar] = _RAND_0[15:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_1[initvar] = _RAND_2[15:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_2[initvar] = _RAND_4[15:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_3[initvar] = _RAND_6[15:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_4[initvar] = _RAND_8[15:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_5[initvar] = _RAND_10[15:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_6[initvar] = _RAND_12[15:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_7[initvar] = _RAND_14[15:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_8[initvar] = _RAND_16[15:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_9[initvar] = _RAND_18[15:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_10[initvar] = _RAND_20[15:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_11[initvar] = _RAND_22[15:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_12[initvar] = _RAND_24[15:0];
  _RAND_26 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_13[initvar] = _RAND_26[15:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_14[initvar] = _RAND_28[15:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_15[initvar] = _RAND_30[15:0];
  _RAND_32 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_16[initvar] = _RAND_32[15:0];
  _RAND_34 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_17[initvar] = _RAND_34[15:0];
  _RAND_36 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_18[initvar] = _RAND_36[15:0];
  _RAND_38 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_19[initvar] = _RAND_38[15:0];
  _RAND_40 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_20[initvar] = _RAND_40[15:0];
  _RAND_42 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_21[initvar] = _RAND_42[15:0];
  _RAND_44 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_22[initvar] = _RAND_44[15:0];
  _RAND_46 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_23[initvar] = _RAND_46[15:0];
  _RAND_48 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_24[initvar] = _RAND_48[15:0];
  _RAND_50 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_25[initvar] = _RAND_50[15:0];
  _RAND_52 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_26[initvar] = _RAND_52[15:0];
  _RAND_54 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_27[initvar] = _RAND_54[15:0];
  _RAND_56 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_28[initvar] = _RAND_56[15:0];
  _RAND_58 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_29[initvar] = _RAND_58[15:0];
  _RAND_60 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_30[initvar] = _RAND_60[15:0];
  _RAND_62 = {1{`RANDOM}};
  for (initvar = 0; initvar < 63; initvar = initvar+1)
    ram_31[initvar] = _RAND_62[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  enq_ptr_value = _RAND_64[5:0];
  _RAND_65 = {1{`RANDOM}};
  deq_ptr_value = _RAND_65[5:0];
  _RAND_66 = {1{`RANDOM}};
  maybe_full = _RAND_66[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SystolicArray(
  input         clock,
  input         reset,
  output        io_control_ready,
  input         io_control_valid,
  input         io_control_bits_load,
  input         io_control_bits_zeroes,
  output        io_input_ready,
  input         io_input_valid,
  input  [15:0] io_input_bits_0,
  input  [15:0] io_input_bits_1,
  input  [15:0] io_input_bits_2,
  input  [15:0] io_input_bits_3,
  input  [15:0] io_input_bits_4,
  input  [15:0] io_input_bits_5,
  input  [15:0] io_input_bits_6,
  input  [15:0] io_input_bits_7,
  input  [15:0] io_input_bits_8,
  input  [15:0] io_input_bits_9,
  input  [15:0] io_input_bits_10,
  input  [15:0] io_input_bits_11,
  input  [15:0] io_input_bits_12,
  input  [15:0] io_input_bits_13,
  input  [15:0] io_input_bits_14,
  input  [15:0] io_input_bits_15,
  input  [15:0] io_input_bits_16,
  input  [15:0] io_input_bits_17,
  input  [15:0] io_input_bits_18,
  input  [15:0] io_input_bits_19,
  input  [15:0] io_input_bits_20,
  input  [15:0] io_input_bits_21,
  input  [15:0] io_input_bits_22,
  input  [15:0] io_input_bits_23,
  input  [15:0] io_input_bits_24,
  input  [15:0] io_input_bits_25,
  input  [15:0] io_input_bits_26,
  input  [15:0] io_input_bits_27,
  input  [15:0] io_input_bits_28,
  input  [15:0] io_input_bits_29,
  input  [15:0] io_input_bits_30,
  input  [15:0] io_input_bits_31,
  output        io_weight_ready,
  input         io_weight_valid,
  input  [15:0] io_weight_bits_0,
  input  [15:0] io_weight_bits_1,
  input  [15:0] io_weight_bits_2,
  input  [15:0] io_weight_bits_3,
  input  [15:0] io_weight_bits_4,
  input  [15:0] io_weight_bits_5,
  input  [15:0] io_weight_bits_6,
  input  [15:0] io_weight_bits_7,
  input  [15:0] io_weight_bits_8,
  input  [15:0] io_weight_bits_9,
  input  [15:0] io_weight_bits_10,
  input  [15:0] io_weight_bits_11,
  input  [15:0] io_weight_bits_12,
  input  [15:0] io_weight_bits_13,
  input  [15:0] io_weight_bits_14,
  input  [15:0] io_weight_bits_15,
  input  [15:0] io_weight_bits_16,
  input  [15:0] io_weight_bits_17,
  input  [15:0] io_weight_bits_18,
  input  [15:0] io_weight_bits_19,
  input  [15:0] io_weight_bits_20,
  input  [15:0] io_weight_bits_21,
  input  [15:0] io_weight_bits_22,
  input  [15:0] io_weight_bits_23,
  input  [15:0] io_weight_bits_24,
  input  [15:0] io_weight_bits_25,
  input  [15:0] io_weight_bits_26,
  input  [15:0] io_weight_bits_27,
  input  [15:0] io_weight_bits_28,
  input  [15:0] io_weight_bits_29,
  input  [15:0] io_weight_bits_30,
  input  [15:0] io_weight_bits_31,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_0,
  output [15:0] io_output_bits_1,
  output [15:0] io_output_bits_2,
  output [15:0] io_output_bits_3,
  output [15:0] io_output_bits_4,
  output [15:0] io_output_bits_5,
  output [15:0] io_output_bits_6,
  output [15:0] io_output_bits_7,
  output [15:0] io_output_bits_8,
  output [15:0] io_output_bits_9,
  output [15:0] io_output_bits_10,
  output [15:0] io_output_bits_11,
  output [15:0] io_output_bits_12,
  output [15:0] io_output_bits_13,
  output [15:0] io_output_bits_14,
  output [15:0] io_output_bits_15,
  output [15:0] io_output_bits_16,
  output [15:0] io_output_bits_17,
  output [15:0] io_output_bits_18,
  output [15:0] io_output_bits_19,
  output [15:0] io_output_bits_20,
  output [15:0] io_output_bits_21,
  output [15:0] io_output_bits_22,
  output [15:0] io_output_bits_23,
  output [15:0] io_output_bits_24,
  output [15:0] io_output_bits_25,
  output [15:0] io_output_bits_26,
  output [15:0] io_output_bits_27,
  output [15:0] io_output_bits_28,
  output [15:0] io_output_bits_29,
  output [15:0] io_output_bits_30,
  output [15:0] io_output_bits_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  wire  array_clock; // @[SystolicArray.scala 40:37]
  wire  array_reset; // @[SystolicArray.scala 40:37]
  wire  array_io_load; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_0; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_1; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_2; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_3; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_4; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_5; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_6; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_7; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_8; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_9; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_10; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_11; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_12; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_13; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_14; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_15; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_16; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_17; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_18; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_19; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_20; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_21; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_22; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_23; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_24; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_25; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_26; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_27; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_28; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_29; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_30; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_input_31; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_0; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_1; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_2; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_3; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_4; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_5; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_6; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_7; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_8; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_9; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_10; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_11; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_12; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_13; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_14; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_15; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_16; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_17; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_18; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_19; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_20; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_21; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_22; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_23; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_24; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_25; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_26; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_27; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_28; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_29; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_30; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_weight_31; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_0; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_1; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_2; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_3; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_4; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_5; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_6; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_7; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_8; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_9; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_10; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_11; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_12; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_13; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_14; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_15; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_16; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_17; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_18; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_19; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_20; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_21; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_22; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_23; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_24; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_25; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_26; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_27; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_28; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_29; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_30; // @[SystolicArray.scala 40:37]
  wire [15:0] array_io_output_31; // @[SystolicArray.scala 40:37]
  wire  output__clock; // @[SystolicArray.scala 45:22]
  wire  output__reset; // @[SystolicArray.scala 45:22]
  wire  output__io_enq_ready; // @[SystolicArray.scala 45:22]
  wire  output__io_enq_valid; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_0; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_1; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_2; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_3; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_4; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_5; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_6; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_7; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_8; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_9; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_10; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_11; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_12; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_13; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_14; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_15; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_16; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_17; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_18; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_19; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_20; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_21; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_22; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_23; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_24; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_25; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_26; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_27; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_28; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_29; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_30; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_enq_bits_31; // @[SystolicArray.scala 45:22]
  wire  output__io_deq_ready; // @[SystolicArray.scala 45:22]
  wire  output__io_deq_valid; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_0; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_1; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_2; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_3; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_4; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_5; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_6; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_7; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_8; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_9; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_10; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_11; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_12; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_13; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_14; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_15; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_16; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_17; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_18; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_19; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_20; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_21; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_22; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_23; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_24; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_25; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_26; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_27; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_28; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_29; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_30; // @[SystolicArray.scala 45:22]
  wire [15:0] output__io_deq_bits_31; // @[SystolicArray.scala 45:22]
  wire  _runInput_T = ~io_control_bits_load; // @[SystolicArray.scala 62:36]
  wire  _runInput_T_1 = io_control_valid & ~io_control_bits_load; // @[SystolicArray.scala 62:33]
  wire  _runInput_T_2 = ~io_control_bits_zeroes; // @[SystolicArray.scala 62:58]
  wire  runInput = io_control_valid & ~io_control_bits_load & ~io_control_bits_zeroes; // @[SystolicArray.scala 62:55]
  wire  runZeroes = _runInput_T_1 & io_control_bits_zeroes; // @[SystolicArray.scala 63:55]
  wire  _loadWeight_T = io_control_valid & io_control_bits_load; // @[SystolicArray.scala 65:19]
  wire  loadWeight = io_control_valid & io_control_bits_load & _runInput_T_2; // @[SystolicArray.scala 65:40]
  wire  loadZeroes = _loadWeight_T & io_control_bits_zeroes; // @[SystolicArray.scala 66:55]
  wire  running = (runInput & io_input_valid & io_input_ready | runZeroes) & output__io_deq_ready; // @[SystolicArray.scala 69:61]
  wire  loading = loadWeight & io_weight_valid & io_weight_ready | loadZeroes; // @[SystolicArray.scala 70:62]
  reg [5:0] arrayPropagationCountdown; // @[SystolicArray.scala 74:42]
  wire [5:0] _arrayPropagationCountdown_T_1 = arrayPropagationCountdown - 6'h1; // @[SystolicArray.scala 81:62]
  wire  inputDone = arrayPropagationCountdown == 6'h0; // @[SystolicArray.scala 87:45]
  wire  _io_control_ready_T_6 = io_control_bits_load & (io_control_bits_zeroes | io_weight_valid) & inputDone; // @[SystolicArray.scala 103:65]
  reg  output_io_enq_valid_sr_0; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_1; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_2; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_3; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_4; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_5; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_6; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_7; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_8; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_9; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_10; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_11; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_12; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_13; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_14; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_15; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_16; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_17; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_18; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_19; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_20; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_21; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_22; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_23; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_24; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_25; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_26; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_27; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_28; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_29; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_30; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_31; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_32; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_33; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_34; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_35; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_36; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_37; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_38; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_39; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_40; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_41; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_42; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_43; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_44; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_45; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_46; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_47; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_48; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_49; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_50; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_51; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_52; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_53; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_54; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_55; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_56; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_57; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_58; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_59; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_60; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_61; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_62; // @[ShiftRegister.scala 10:22]
  InnerSystolicArray array ( // @[SystolicArray.scala 40:37]
    .clock(array_clock),
    .reset(array_reset),
    .io_load(array_io_load),
    .io_input_0(array_io_input_0),
    .io_input_1(array_io_input_1),
    .io_input_2(array_io_input_2),
    .io_input_3(array_io_input_3),
    .io_input_4(array_io_input_4),
    .io_input_5(array_io_input_5),
    .io_input_6(array_io_input_6),
    .io_input_7(array_io_input_7),
    .io_input_8(array_io_input_8),
    .io_input_9(array_io_input_9),
    .io_input_10(array_io_input_10),
    .io_input_11(array_io_input_11),
    .io_input_12(array_io_input_12),
    .io_input_13(array_io_input_13),
    .io_input_14(array_io_input_14),
    .io_input_15(array_io_input_15),
    .io_input_16(array_io_input_16),
    .io_input_17(array_io_input_17),
    .io_input_18(array_io_input_18),
    .io_input_19(array_io_input_19),
    .io_input_20(array_io_input_20),
    .io_input_21(array_io_input_21),
    .io_input_22(array_io_input_22),
    .io_input_23(array_io_input_23),
    .io_input_24(array_io_input_24),
    .io_input_25(array_io_input_25),
    .io_input_26(array_io_input_26),
    .io_input_27(array_io_input_27),
    .io_input_28(array_io_input_28),
    .io_input_29(array_io_input_29),
    .io_input_30(array_io_input_30),
    .io_input_31(array_io_input_31),
    .io_weight_0(array_io_weight_0),
    .io_weight_1(array_io_weight_1),
    .io_weight_2(array_io_weight_2),
    .io_weight_3(array_io_weight_3),
    .io_weight_4(array_io_weight_4),
    .io_weight_5(array_io_weight_5),
    .io_weight_6(array_io_weight_6),
    .io_weight_7(array_io_weight_7),
    .io_weight_8(array_io_weight_8),
    .io_weight_9(array_io_weight_9),
    .io_weight_10(array_io_weight_10),
    .io_weight_11(array_io_weight_11),
    .io_weight_12(array_io_weight_12),
    .io_weight_13(array_io_weight_13),
    .io_weight_14(array_io_weight_14),
    .io_weight_15(array_io_weight_15),
    .io_weight_16(array_io_weight_16),
    .io_weight_17(array_io_weight_17),
    .io_weight_18(array_io_weight_18),
    .io_weight_19(array_io_weight_19),
    .io_weight_20(array_io_weight_20),
    .io_weight_21(array_io_weight_21),
    .io_weight_22(array_io_weight_22),
    .io_weight_23(array_io_weight_23),
    .io_weight_24(array_io_weight_24),
    .io_weight_25(array_io_weight_25),
    .io_weight_26(array_io_weight_26),
    .io_weight_27(array_io_weight_27),
    .io_weight_28(array_io_weight_28),
    .io_weight_29(array_io_weight_29),
    .io_weight_30(array_io_weight_30),
    .io_weight_31(array_io_weight_31),
    .io_output_0(array_io_output_0),
    .io_output_1(array_io_output_1),
    .io_output_2(array_io_output_2),
    .io_output_3(array_io_output_3),
    .io_output_4(array_io_output_4),
    .io_output_5(array_io_output_5),
    .io_output_6(array_io_output_6),
    .io_output_7(array_io_output_7),
    .io_output_8(array_io_output_8),
    .io_output_9(array_io_output_9),
    .io_output_10(array_io_output_10),
    .io_output_11(array_io_output_11),
    .io_output_12(array_io_output_12),
    .io_output_13(array_io_output_13),
    .io_output_14(array_io_output_14),
    .io_output_15(array_io_output_15),
    .io_output_16(array_io_output_16),
    .io_output_17(array_io_output_17),
    .io_output_18(array_io_output_18),
    .io_output_19(array_io_output_19),
    .io_output_20(array_io_output_20),
    .io_output_21(array_io_output_21),
    .io_output_22(array_io_output_22),
    .io_output_23(array_io_output_23),
    .io_output_24(array_io_output_24),
    .io_output_25(array_io_output_25),
    .io_output_26(array_io_output_26),
    .io_output_27(array_io_output_27),
    .io_output_28(array_io_output_28),
    .io_output_29(array_io_output_29),
    .io_output_30(array_io_output_30),
    .io_output_31(array_io_output_31)
  );
  Queue_8 output_ ( // @[SystolicArray.scala 45:22]
    .clock(output__clock),
    .reset(output__reset),
    .io_enq_ready(output__io_enq_ready),
    .io_enq_valid(output__io_enq_valid),
    .io_enq_bits_0(output__io_enq_bits_0),
    .io_enq_bits_1(output__io_enq_bits_1),
    .io_enq_bits_2(output__io_enq_bits_2),
    .io_enq_bits_3(output__io_enq_bits_3),
    .io_enq_bits_4(output__io_enq_bits_4),
    .io_enq_bits_5(output__io_enq_bits_5),
    .io_enq_bits_6(output__io_enq_bits_6),
    .io_enq_bits_7(output__io_enq_bits_7),
    .io_enq_bits_8(output__io_enq_bits_8),
    .io_enq_bits_9(output__io_enq_bits_9),
    .io_enq_bits_10(output__io_enq_bits_10),
    .io_enq_bits_11(output__io_enq_bits_11),
    .io_enq_bits_12(output__io_enq_bits_12),
    .io_enq_bits_13(output__io_enq_bits_13),
    .io_enq_bits_14(output__io_enq_bits_14),
    .io_enq_bits_15(output__io_enq_bits_15),
    .io_enq_bits_16(output__io_enq_bits_16),
    .io_enq_bits_17(output__io_enq_bits_17),
    .io_enq_bits_18(output__io_enq_bits_18),
    .io_enq_bits_19(output__io_enq_bits_19),
    .io_enq_bits_20(output__io_enq_bits_20),
    .io_enq_bits_21(output__io_enq_bits_21),
    .io_enq_bits_22(output__io_enq_bits_22),
    .io_enq_bits_23(output__io_enq_bits_23),
    .io_enq_bits_24(output__io_enq_bits_24),
    .io_enq_bits_25(output__io_enq_bits_25),
    .io_enq_bits_26(output__io_enq_bits_26),
    .io_enq_bits_27(output__io_enq_bits_27),
    .io_enq_bits_28(output__io_enq_bits_28),
    .io_enq_bits_29(output__io_enq_bits_29),
    .io_enq_bits_30(output__io_enq_bits_30),
    .io_enq_bits_31(output__io_enq_bits_31),
    .io_deq_ready(output__io_deq_ready),
    .io_deq_valid(output__io_deq_valid),
    .io_deq_bits_0(output__io_deq_bits_0),
    .io_deq_bits_1(output__io_deq_bits_1),
    .io_deq_bits_2(output__io_deq_bits_2),
    .io_deq_bits_3(output__io_deq_bits_3),
    .io_deq_bits_4(output__io_deq_bits_4),
    .io_deq_bits_5(output__io_deq_bits_5),
    .io_deq_bits_6(output__io_deq_bits_6),
    .io_deq_bits_7(output__io_deq_bits_7),
    .io_deq_bits_8(output__io_deq_bits_8),
    .io_deq_bits_9(output__io_deq_bits_9),
    .io_deq_bits_10(output__io_deq_bits_10),
    .io_deq_bits_11(output__io_deq_bits_11),
    .io_deq_bits_12(output__io_deq_bits_12),
    .io_deq_bits_13(output__io_deq_bits_13),
    .io_deq_bits_14(output__io_deq_bits_14),
    .io_deq_bits_15(output__io_deq_bits_15),
    .io_deq_bits_16(output__io_deq_bits_16),
    .io_deq_bits_17(output__io_deq_bits_17),
    .io_deq_bits_18(output__io_deq_bits_18),
    .io_deq_bits_19(output__io_deq_bits_19),
    .io_deq_bits_20(output__io_deq_bits_20),
    .io_deq_bits_21(output__io_deq_bits_21),
    .io_deq_bits_22(output__io_deq_bits_22),
    .io_deq_bits_23(output__io_deq_bits_23),
    .io_deq_bits_24(output__io_deq_bits_24),
    .io_deq_bits_25(output__io_deq_bits_25),
    .io_deq_bits_26(output__io_deq_bits_26),
    .io_deq_bits_27(output__io_deq_bits_27),
    .io_deq_bits_28(output__io_deq_bits_28),
    .io_deq_bits_29(output__io_deq_bits_29),
    .io_deq_bits_30(output__io_deq_bits_30),
    .io_deq_bits_31(output__io_deq_bits_31)
  );
  assign io_control_ready = _runInput_T & (io_control_bits_zeroes | io_input_valid) & output__io_deq_ready |
    _io_control_ready_T_6; // @[SystolicArray.scala 102:104]
  assign io_input_ready = runInput & output__io_deq_ready; // @[SystolicArray.scala 100:27]
  assign io_weight_ready = loadWeight & inputDone; // @[SystolicArray.scala 101:30]
  assign io_output_valid = output__io_deq_valid; // @[SystolicArray.scala 98:13]
  assign io_output_bits_0 = output__io_deq_bits_0; // @[SystolicArray.scala 98:13]
  assign io_output_bits_1 = output__io_deq_bits_1; // @[SystolicArray.scala 98:13]
  assign io_output_bits_2 = output__io_deq_bits_2; // @[SystolicArray.scala 98:13]
  assign io_output_bits_3 = output__io_deq_bits_3; // @[SystolicArray.scala 98:13]
  assign io_output_bits_4 = output__io_deq_bits_4; // @[SystolicArray.scala 98:13]
  assign io_output_bits_5 = output__io_deq_bits_5; // @[SystolicArray.scala 98:13]
  assign io_output_bits_6 = output__io_deq_bits_6; // @[SystolicArray.scala 98:13]
  assign io_output_bits_7 = output__io_deq_bits_7; // @[SystolicArray.scala 98:13]
  assign io_output_bits_8 = output__io_deq_bits_8; // @[SystolicArray.scala 98:13]
  assign io_output_bits_9 = output__io_deq_bits_9; // @[SystolicArray.scala 98:13]
  assign io_output_bits_10 = output__io_deq_bits_10; // @[SystolicArray.scala 98:13]
  assign io_output_bits_11 = output__io_deq_bits_11; // @[SystolicArray.scala 98:13]
  assign io_output_bits_12 = output__io_deq_bits_12; // @[SystolicArray.scala 98:13]
  assign io_output_bits_13 = output__io_deq_bits_13; // @[SystolicArray.scala 98:13]
  assign io_output_bits_14 = output__io_deq_bits_14; // @[SystolicArray.scala 98:13]
  assign io_output_bits_15 = output__io_deq_bits_15; // @[SystolicArray.scala 98:13]
  assign io_output_bits_16 = output__io_deq_bits_16; // @[SystolicArray.scala 98:13]
  assign io_output_bits_17 = output__io_deq_bits_17; // @[SystolicArray.scala 98:13]
  assign io_output_bits_18 = output__io_deq_bits_18; // @[SystolicArray.scala 98:13]
  assign io_output_bits_19 = output__io_deq_bits_19; // @[SystolicArray.scala 98:13]
  assign io_output_bits_20 = output__io_deq_bits_20; // @[SystolicArray.scala 98:13]
  assign io_output_bits_21 = output__io_deq_bits_21; // @[SystolicArray.scala 98:13]
  assign io_output_bits_22 = output__io_deq_bits_22; // @[SystolicArray.scala 98:13]
  assign io_output_bits_23 = output__io_deq_bits_23; // @[SystolicArray.scala 98:13]
  assign io_output_bits_24 = output__io_deq_bits_24; // @[SystolicArray.scala 98:13]
  assign io_output_bits_25 = output__io_deq_bits_25; // @[SystolicArray.scala 98:13]
  assign io_output_bits_26 = output__io_deq_bits_26; // @[SystolicArray.scala 98:13]
  assign io_output_bits_27 = output__io_deq_bits_27; // @[SystolicArray.scala 98:13]
  assign io_output_bits_28 = output__io_deq_bits_28; // @[SystolicArray.scala 98:13]
  assign io_output_bits_29 = output__io_deq_bits_29; // @[SystolicArray.scala 98:13]
  assign io_output_bits_30 = output__io_deq_bits_30; // @[SystolicArray.scala 98:13]
  assign io_output_bits_31 = output__io_deq_bits_31; // @[SystolicArray.scala 98:13]
  assign array_clock = clock;
  assign array_reset = reset;
  assign array_io_load = inputDone & loading; // @[SystolicArray.scala 89:30]
  assign array_io_input_0 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_0); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_1 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_1); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_2 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_2); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_3 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_3); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_4 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_4); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_5 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_5); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_6 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_6); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_7 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_7); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_8 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_8); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_9 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_9); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_10 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_10); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_11 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_11); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_12 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_12); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_13 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_13); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_14 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_14); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_15 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_15); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_16 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_16); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_17 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_17); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_18 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_18); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_19 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_19); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_20 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_20); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_21 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_21); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_22 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_22); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_23 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_23); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_24 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_24); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_25 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_25); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_26 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_26); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_27 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_27); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_28 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_28); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_29 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_29); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_30 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_30); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_input_31 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_input_bits_31); // @[SystolicArray.scala 90:29 91:20 94:20]
  assign array_io_weight_0 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_0); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_1 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_1); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_2 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_2); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_3 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_3); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_4 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_4); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_5 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_5); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_6 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_6); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_7 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_7); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_8 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_8); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_9 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_9); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_10 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_10); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_11 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_11); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_12 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_12); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_13 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_13); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_14 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_14); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_15 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_15); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_16 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_16); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_17 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_17); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_18 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_18); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_19 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_19); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_20 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_20); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_21 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_21); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_22 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_22); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_23 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_23); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_24 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_24); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_25 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_25); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_26 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_26); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_27 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_27); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_28 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_28); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_29 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_29); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_30 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_30); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign array_io_weight_31 = io_control_bits_zeroes ? $signed(16'sh0) : $signed(io_weight_bits_31); // @[SystolicArray.scala 90:29 92:21 95:21]
  assign output__clock = clock;
  assign output__reset = reset;
  assign output__io_enq_valid = output_io_enq_valid_sr_62; // @[SystolicArray.scala 106:23]
  assign output__io_enq_bits_0 = array_io_output_0; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_1 = array_io_output_1; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_2 = array_io_output_2; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_3 = array_io_output_3; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_4 = array_io_output_4; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_5 = array_io_output_5; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_6 = array_io_output_6; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_7 = array_io_output_7; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_8 = array_io_output_8; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_9 = array_io_output_9; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_10 = array_io_output_10; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_11 = array_io_output_11; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_12 = array_io_output_12; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_13 = array_io_output_13; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_14 = array_io_output_14; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_15 = array_io_output_15; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_16 = array_io_output_16; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_17 = array_io_output_17; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_18 = array_io_output_18; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_19 = array_io_output_19; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_20 = array_io_output_20; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_21 = array_io_output_21; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_22 = array_io_output_22; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_23 = array_io_output_23; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_24 = array_io_output_24; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_25 = array_io_output_25; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_26 = array_io_output_26; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_27 = array_io_output_27; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_28 = array_io_output_28; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_29 = array_io_output_29; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_30 = array_io_output_30; // @[SystolicArray.scala 97:22]
  assign output__io_enq_bits_31 = array_io_output_31; // @[SystolicArray.scala 97:22]
  assign output__io_deq_ready = io_output_ready; // @[SystolicArray.scala 98:13]
  always @(posedge clock) begin
    if (reset) begin // @[SystolicArray.scala 74:42]
      arrayPropagationCountdown <= 6'h0; // @[SystolicArray.scala 74:42]
    end else if (running) begin // @[SystolicArray.scala 77:17]
      arrayPropagationCountdown <= 6'h3f; // @[SystolicArray.scala 78:31]
    end else if (arrayPropagationCountdown > 6'h0) begin // @[SystolicArray.scala 80:43]
      arrayPropagationCountdown <= _arrayPropagationCountdown_T_1; // @[SystolicArray.scala 81:33]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_0 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_0 <= running; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_1 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_1 <= output_io_enq_valid_sr_0; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_2 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_2 <= output_io_enq_valid_sr_1; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_3 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_3 <= output_io_enq_valid_sr_2; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_4 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_4 <= output_io_enq_valid_sr_3; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_5 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_5 <= output_io_enq_valid_sr_4; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_6 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_6 <= output_io_enq_valid_sr_5; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_7 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_7 <= output_io_enq_valid_sr_6; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_8 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_8 <= output_io_enq_valid_sr_7; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_9 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_9 <= output_io_enq_valid_sr_8; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_10 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_10 <= output_io_enq_valid_sr_9; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_11 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_11 <= output_io_enq_valid_sr_10; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_12 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_12 <= output_io_enq_valid_sr_11; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_13 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_13 <= output_io_enq_valid_sr_12; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_14 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_14 <= output_io_enq_valid_sr_13; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_15 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_15 <= output_io_enq_valid_sr_14; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_16 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_16 <= output_io_enq_valid_sr_15; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_17 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_17 <= output_io_enq_valid_sr_16; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_18 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_18 <= output_io_enq_valid_sr_17; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_19 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_19 <= output_io_enq_valid_sr_18; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_20 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_20 <= output_io_enq_valid_sr_19; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_21 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_21 <= output_io_enq_valid_sr_20; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_22 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_22 <= output_io_enq_valid_sr_21; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_23 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_23 <= output_io_enq_valid_sr_22; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_24 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_24 <= output_io_enq_valid_sr_23; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_25 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_25 <= output_io_enq_valid_sr_24; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_26 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_26 <= output_io_enq_valid_sr_25; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_27 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_27 <= output_io_enq_valid_sr_26; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_28 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_28 <= output_io_enq_valid_sr_27; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_29 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_29 <= output_io_enq_valid_sr_28; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_30 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_30 <= output_io_enq_valid_sr_29; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_31 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_31 <= output_io_enq_valid_sr_30; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_32 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_32 <= output_io_enq_valid_sr_31; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_33 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_33 <= output_io_enq_valid_sr_32; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_34 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_34 <= output_io_enq_valid_sr_33; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_35 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_35 <= output_io_enq_valid_sr_34; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_36 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_36 <= output_io_enq_valid_sr_35; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_37 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_37 <= output_io_enq_valid_sr_36; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_38 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_38 <= output_io_enq_valid_sr_37; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_39 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_39 <= output_io_enq_valid_sr_38; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_40 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_40 <= output_io_enq_valid_sr_39; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_41 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_41 <= output_io_enq_valid_sr_40; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_42 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_42 <= output_io_enq_valid_sr_41; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_43 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_43 <= output_io_enq_valid_sr_42; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_44 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_44 <= output_io_enq_valid_sr_43; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_45 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_45 <= output_io_enq_valid_sr_44; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_46 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_46 <= output_io_enq_valid_sr_45; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_47 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_47 <= output_io_enq_valid_sr_46; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_48 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_48 <= output_io_enq_valid_sr_47; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_49 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_49 <= output_io_enq_valid_sr_48; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_50 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_50 <= output_io_enq_valid_sr_49; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_51 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_51 <= output_io_enq_valid_sr_50; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_52 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_52 <= output_io_enq_valid_sr_51; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_53 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_53 <= output_io_enq_valid_sr_52; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_54 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_54 <= output_io_enq_valid_sr_53; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_55 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_55 <= output_io_enq_valid_sr_54; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_56 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_56 <= output_io_enq_valid_sr_55; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_57 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_57 <= output_io_enq_valid_sr_56; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_58 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_58 <= output_io_enq_valid_sr_57; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_59 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_59 <= output_io_enq_valid_sr_58; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_60 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_60 <= output_io_enq_valid_sr_59; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_61 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_61 <= output_io_enq_valid_sr_60; // @[ShiftRegister.scala 13:11]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_62 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_62 <= output_io_enq_valid_sr_61; // @[ShiftRegister.scala 13:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  arrayPropagationCountdown = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  output_io_enq_valid_sr_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  output_io_enq_valid_sr_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  output_io_enq_valid_sr_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  output_io_enq_valid_sr_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  output_io_enq_valid_sr_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  output_io_enq_valid_sr_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  output_io_enq_valid_sr_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  output_io_enq_valid_sr_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  output_io_enq_valid_sr_8 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  output_io_enq_valid_sr_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  output_io_enq_valid_sr_10 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  output_io_enq_valid_sr_11 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  output_io_enq_valid_sr_12 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  output_io_enq_valid_sr_13 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  output_io_enq_valid_sr_14 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  output_io_enq_valid_sr_15 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  output_io_enq_valid_sr_16 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  output_io_enq_valid_sr_17 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  output_io_enq_valid_sr_18 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  output_io_enq_valid_sr_19 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  output_io_enq_valid_sr_20 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  output_io_enq_valid_sr_21 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  output_io_enq_valid_sr_22 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  output_io_enq_valid_sr_23 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  output_io_enq_valid_sr_24 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  output_io_enq_valid_sr_25 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  output_io_enq_valid_sr_26 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  output_io_enq_valid_sr_27 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  output_io_enq_valid_sr_28 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  output_io_enq_valid_sr_29 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  output_io_enq_valid_sr_30 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  output_io_enq_valid_sr_31 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  output_io_enq_valid_sr_32 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  output_io_enq_valid_sr_33 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  output_io_enq_valid_sr_34 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  output_io_enq_valid_sr_35 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  output_io_enq_valid_sr_36 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  output_io_enq_valid_sr_37 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  output_io_enq_valid_sr_38 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  output_io_enq_valid_sr_39 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  output_io_enq_valid_sr_40 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  output_io_enq_valid_sr_41 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  output_io_enq_valid_sr_42 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  output_io_enq_valid_sr_43 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  output_io_enq_valid_sr_44 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  output_io_enq_valid_sr_45 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  output_io_enq_valid_sr_46 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  output_io_enq_valid_sr_47 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  output_io_enq_valid_sr_48 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  output_io_enq_valid_sr_49 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  output_io_enq_valid_sr_50 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  output_io_enq_valid_sr_51 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  output_io_enq_valid_sr_52 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  output_io_enq_valid_sr_53 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  output_io_enq_valid_sr_54 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  output_io_enq_valid_sr_55 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  output_io_enq_valid_sr_56 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  output_io_enq_valid_sr_57 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  output_io_enq_valid_sr_58 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  output_io_enq_valid_sr_59 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  output_io_enq_valid_sr_60 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  output_io_enq_valid_sr_61 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  output_io_enq_valid_sr_62 = _RAND_63[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InnerDualPortMem(
  input         clock,
  input         reset,
  input  [11:0] io_portA_address,
  input         io_portA_read_enable,
  output [15:0] io_portA_read_data_0,
  output [15:0] io_portA_read_data_1,
  output [15:0] io_portA_read_data_2,
  output [15:0] io_portA_read_data_3,
  output [15:0] io_portA_read_data_4,
  output [15:0] io_portA_read_data_5,
  output [15:0] io_portA_read_data_6,
  output [15:0] io_portA_read_data_7,
  output [15:0] io_portA_read_data_8,
  output [15:0] io_portA_read_data_9,
  output [15:0] io_portA_read_data_10,
  output [15:0] io_portA_read_data_11,
  output [15:0] io_portA_read_data_12,
  output [15:0] io_portA_read_data_13,
  output [15:0] io_portA_read_data_14,
  output [15:0] io_portA_read_data_15,
  output [15:0] io_portA_read_data_16,
  output [15:0] io_portA_read_data_17,
  output [15:0] io_portA_read_data_18,
  output [15:0] io_portA_read_data_19,
  output [15:0] io_portA_read_data_20,
  output [15:0] io_portA_read_data_21,
  output [15:0] io_portA_read_data_22,
  output [15:0] io_portA_read_data_23,
  output [15:0] io_portA_read_data_24,
  output [15:0] io_portA_read_data_25,
  output [15:0] io_portA_read_data_26,
  output [15:0] io_portA_read_data_27,
  output [15:0] io_portA_read_data_28,
  output [15:0] io_portA_read_data_29,
  output [15:0] io_portA_read_data_30,
  output [15:0] io_portA_read_data_31,
  input         io_portA_write_enable,
  input  [15:0] io_portA_write_data_0,
  input  [15:0] io_portA_write_data_1,
  input  [15:0] io_portA_write_data_2,
  input  [15:0] io_portA_write_data_3,
  input  [15:0] io_portA_write_data_4,
  input  [15:0] io_portA_write_data_5,
  input  [15:0] io_portA_write_data_6,
  input  [15:0] io_portA_write_data_7,
  input  [15:0] io_portA_write_data_8,
  input  [15:0] io_portA_write_data_9,
  input  [15:0] io_portA_write_data_10,
  input  [15:0] io_portA_write_data_11,
  input  [15:0] io_portA_write_data_12,
  input  [15:0] io_portA_write_data_13,
  input  [15:0] io_portA_write_data_14,
  input  [15:0] io_portA_write_data_15,
  input  [15:0] io_portA_write_data_16,
  input  [15:0] io_portA_write_data_17,
  input  [15:0] io_portA_write_data_18,
  input  [15:0] io_portA_write_data_19,
  input  [15:0] io_portA_write_data_20,
  input  [15:0] io_portA_write_data_21,
  input  [15:0] io_portA_write_data_22,
  input  [15:0] io_portA_write_data_23,
  input  [15:0] io_portA_write_data_24,
  input  [15:0] io_portA_write_data_25,
  input  [15:0] io_portA_write_data_26,
  input  [15:0] io_portA_write_data_27,
  input  [15:0] io_portA_write_data_28,
  input  [15:0] io_portA_write_data_29,
  input  [15:0] io_portA_write_data_30,
  input  [15:0] io_portA_write_data_31,
  input  [11:0] io_portB_address,
  input         io_portB_read_enable,
  output [15:0] io_portB_read_data_0,
  output [15:0] io_portB_read_data_1,
  output [15:0] io_portB_read_data_2,
  output [15:0] io_portB_read_data_3,
  output [15:0] io_portB_read_data_4,
  output [15:0] io_portB_read_data_5,
  output [15:0] io_portB_read_data_6,
  output [15:0] io_portB_read_data_7,
  output [15:0] io_portB_read_data_8,
  output [15:0] io_portB_read_data_9,
  output [15:0] io_portB_read_data_10,
  output [15:0] io_portB_read_data_11,
  output [15:0] io_portB_read_data_12,
  output [15:0] io_portB_read_data_13,
  output [15:0] io_portB_read_data_14,
  output [15:0] io_portB_read_data_15,
  output [15:0] io_portB_read_data_16,
  output [15:0] io_portB_read_data_17,
  output [15:0] io_portB_read_data_18,
  output [15:0] io_portB_read_data_19,
  output [15:0] io_portB_read_data_20,
  output [15:0] io_portB_read_data_21,
  output [15:0] io_portB_read_data_22,
  output [15:0] io_portB_read_data_23,
  output [15:0] io_portB_read_data_24,
  output [15:0] io_portB_read_data_25,
  output [15:0] io_portB_read_data_26,
  output [15:0] io_portB_read_data_27,
  output [15:0] io_portB_read_data_28,
  output [15:0] io_portB_read_data_29,
  output [15:0] io_portB_read_data_30,
  output [15:0] io_portB_read_data_31
);
  wire  mem_clka; // @[DualPortMem.scala 173:25]
  wire  mem_wea; // @[DualPortMem.scala 173:25]
  wire  mem_ena; // @[DualPortMem.scala 173:25]
  wire [11:0] mem_addra; // @[DualPortMem.scala 173:25]
  wire [511:0] mem_dia; // @[DualPortMem.scala 173:25]
  wire [511:0] mem_doa; // @[DualPortMem.scala 173:25]
  wire  mem_clkb; // @[DualPortMem.scala 173:25]
  wire  mem_web; // @[DualPortMem.scala 173:25]
  wire  mem_enb; // @[DualPortMem.scala 173:25]
  wire [11:0] mem_addrb; // @[DualPortMem.scala 173:25]
  wire [511:0] mem_dib; // @[DualPortMem.scala 173:25]
  wire [511:0] mem_dob; // @[DualPortMem.scala 173:25]
  wire [511:0] _io_portA_read_data_WIRE_1 = mem_doa;
  wire [127:0] mem_io_dia_lo_lo = {io_portA_write_data_7,io_portA_write_data_6,io_portA_write_data_5,
    io_portA_write_data_4,io_portA_write_data_3,io_portA_write_data_2,io_portA_write_data_1,io_portA_write_data_0}; // @[DualPortMem.scala 180:51]
  wire [255:0] mem_io_dia_lo = {io_portA_write_data_15,io_portA_write_data_14,io_portA_write_data_13,
    io_portA_write_data_12,io_portA_write_data_11,io_portA_write_data_10,io_portA_write_data_9,io_portA_write_data_8,
    mem_io_dia_lo_lo}; // @[DualPortMem.scala 180:51]
  wire [127:0] mem_io_dia_hi_lo = {io_portA_write_data_23,io_portA_write_data_22,io_portA_write_data_21,
    io_portA_write_data_20,io_portA_write_data_19,io_portA_write_data_18,io_portA_write_data_17,io_portA_write_data_16}; // @[DualPortMem.scala 180:51]
  wire [255:0] mem_io_dia_hi = {io_portA_write_data_31,io_portA_write_data_30,io_portA_write_data_29,
    io_portA_write_data_28,io_portA_write_data_27,io_portA_write_data_26,io_portA_write_data_25,io_portA_write_data_24,
    mem_io_dia_hi_lo}; // @[DualPortMem.scala 180:51]
  wire [511:0] _io_portB_read_data_WIRE_1 = mem_dob;
  bram_dp_512x4096 mem ( // @[DualPortMem.scala 173:25]
    .clka(mem_clka),
    .wea(mem_wea),
    .ena(mem_ena),
    .addra(mem_addra),
    .dia(mem_dia),
    .doa(mem_doa),
    .clkb(mem_clkb),
    .web(mem_web),
    .enb(mem_enb),
    .addrb(mem_addrb),
    .dib(mem_dib),
    .dob(mem_dob)
  );
  assign io_portA_read_data_0 = _io_portA_read_data_WIRE_1[15:0]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_1 = _io_portA_read_data_WIRE_1[31:16]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_2 = _io_portA_read_data_WIRE_1[47:32]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_3 = _io_portA_read_data_WIRE_1[63:48]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_4 = _io_portA_read_data_WIRE_1[79:64]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_5 = _io_portA_read_data_WIRE_1[95:80]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_6 = _io_portA_read_data_WIRE_1[111:96]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_7 = _io_portA_read_data_WIRE_1[127:112]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_8 = _io_portA_read_data_WIRE_1[143:128]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_9 = _io_portA_read_data_WIRE_1[159:144]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_10 = _io_portA_read_data_WIRE_1[175:160]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_11 = _io_portA_read_data_WIRE_1[191:176]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_12 = _io_portA_read_data_WIRE_1[207:192]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_13 = _io_portA_read_data_WIRE_1[223:208]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_14 = _io_portA_read_data_WIRE_1[239:224]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_15 = _io_portA_read_data_WIRE_1[255:240]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_16 = _io_portA_read_data_WIRE_1[271:256]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_17 = _io_portA_read_data_WIRE_1[287:272]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_18 = _io_portA_read_data_WIRE_1[303:288]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_19 = _io_portA_read_data_WIRE_1[319:304]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_20 = _io_portA_read_data_WIRE_1[335:320]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_21 = _io_portA_read_data_WIRE_1[351:336]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_22 = _io_portA_read_data_WIRE_1[367:352]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_23 = _io_portA_read_data_WIRE_1[383:368]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_24 = _io_portA_read_data_WIRE_1[399:384]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_25 = _io_portA_read_data_WIRE_1[415:400]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_26 = _io_portA_read_data_WIRE_1[431:416]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_27 = _io_portA_read_data_WIRE_1[447:432]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_28 = _io_portA_read_data_WIRE_1[463:448]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_29 = _io_portA_read_data_WIRE_1[479:464]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_30 = _io_portA_read_data_WIRE_1[495:480]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_31 = _io_portA_read_data_WIRE_1[511:496]; // @[DualPortMem.scala 178:50]
  assign io_portB_read_data_0 = _io_portB_read_data_WIRE_1[15:0]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_1 = _io_portB_read_data_WIRE_1[31:16]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_2 = _io_portB_read_data_WIRE_1[47:32]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_3 = _io_portB_read_data_WIRE_1[63:48]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_4 = _io_portB_read_data_WIRE_1[79:64]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_5 = _io_portB_read_data_WIRE_1[95:80]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_6 = _io_portB_read_data_WIRE_1[111:96]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_7 = _io_portB_read_data_WIRE_1[127:112]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_8 = _io_portB_read_data_WIRE_1[143:128]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_9 = _io_portB_read_data_WIRE_1[159:144]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_10 = _io_portB_read_data_WIRE_1[175:160]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_11 = _io_portB_read_data_WIRE_1[191:176]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_12 = _io_portB_read_data_WIRE_1[207:192]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_13 = _io_portB_read_data_WIRE_1[223:208]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_14 = _io_portB_read_data_WIRE_1[239:224]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_15 = _io_portB_read_data_WIRE_1[255:240]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_16 = _io_portB_read_data_WIRE_1[271:256]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_17 = _io_portB_read_data_WIRE_1[287:272]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_18 = _io_portB_read_data_WIRE_1[303:288]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_19 = _io_portB_read_data_WIRE_1[319:304]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_20 = _io_portB_read_data_WIRE_1[335:320]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_21 = _io_portB_read_data_WIRE_1[351:336]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_22 = _io_portB_read_data_WIRE_1[367:352]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_23 = _io_portB_read_data_WIRE_1[383:368]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_24 = _io_portB_read_data_WIRE_1[399:384]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_25 = _io_portB_read_data_WIRE_1[415:400]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_26 = _io_portB_read_data_WIRE_1[431:416]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_27 = _io_portB_read_data_WIRE_1[447:432]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_28 = _io_portB_read_data_WIRE_1[463:448]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_29 = _io_portB_read_data_WIRE_1[479:464]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_30 = _io_portB_read_data_WIRE_1[495:480]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_31 = _io_portB_read_data_WIRE_1[511:496]; // @[DualPortMem.scala 185:50]
  assign mem_clka = clock; // @[DualPortMem.scala 175:30]
  assign mem_wea = io_portA_write_enable; // @[DualPortMem.scala 179:20]
  assign mem_ena = ~reset; // @[DualPortMem.scala 176:23]
  assign mem_addra = io_portA_address; // @[DualPortMem.scala 177:22]
  assign mem_dia = {mem_io_dia_hi,mem_io_dia_lo}; // @[DualPortMem.scala 180:51]
  assign mem_clkb = clock; // @[DualPortMem.scala 182:30]
  assign mem_web = 1'h0; // @[DualPortMem.scala 186:20]
  assign mem_enb = ~reset; // @[DualPortMem.scala 183:23]
  assign mem_addrb = io_portB_address; // @[DualPortMem.scala 184:22]
  assign mem_dib = 512'h0; // @[DualPortMem.scala 187:51]
endmodule
module Queue_10(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_0,
  input  [15:0] io_enq_bits_1,
  input  [15:0] io_enq_bits_2,
  input  [15:0] io_enq_bits_3,
  input  [15:0] io_enq_bits_4,
  input  [15:0] io_enq_bits_5,
  input  [15:0] io_enq_bits_6,
  input  [15:0] io_enq_bits_7,
  input  [15:0] io_enq_bits_8,
  input  [15:0] io_enq_bits_9,
  input  [15:0] io_enq_bits_10,
  input  [15:0] io_enq_bits_11,
  input  [15:0] io_enq_bits_12,
  input  [15:0] io_enq_bits_13,
  input  [15:0] io_enq_bits_14,
  input  [15:0] io_enq_bits_15,
  input  [15:0] io_enq_bits_16,
  input  [15:0] io_enq_bits_17,
  input  [15:0] io_enq_bits_18,
  input  [15:0] io_enq_bits_19,
  input  [15:0] io_enq_bits_20,
  input  [15:0] io_enq_bits_21,
  input  [15:0] io_enq_bits_22,
  input  [15:0] io_enq_bits_23,
  input  [15:0] io_enq_bits_24,
  input  [15:0] io_enq_bits_25,
  input  [15:0] io_enq_bits_26,
  input  [15:0] io_enq_bits_27,
  input  [15:0] io_enq_bits_28,
  input  [15:0] io_enq_bits_29,
  input  [15:0] io_enq_bits_30,
  input  [15:0] io_enq_bits_31,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_0,
  output [15:0] io_deq_bits_1,
  output [15:0] io_deq_bits_2,
  output [15:0] io_deq_bits_3,
  output [15:0] io_deq_bits_4,
  output [15:0] io_deq_bits_5,
  output [15:0] io_deq_bits_6,
  output [15:0] io_deq_bits_7,
  output [15:0] io_deq_bits_8,
  output [15:0] io_deq_bits_9,
  output [15:0] io_deq_bits_10,
  output [15:0] io_deq_bits_11,
  output [15:0] io_deq_bits_12,
  output [15:0] io_deq_bits_13,
  output [15:0] io_deq_bits_14,
  output [15:0] io_deq_bits_15,
  output [15:0] io_deq_bits_16,
  output [15:0] io_deq_bits_17,
  output [15:0] io_deq_bits_18,
  output [15:0] io_deq_bits_19,
  output [15:0] io_deq_bits_20,
  output [15:0] io_deq_bits_21,
  output [15:0] io_deq_bits_22,
  output [15:0] io_deq_bits_23,
  output [15:0] io_deq_bits_24,
  output [15:0] io_deq_bits_25,
  output [15:0] io_deq_bits_26,
  output [15:0] io_deq_bits_27,
  output [15:0] io_deq_bits_28,
  output [15:0] io_deq_bits_29,
  output [15:0] io_deq_bits_30,
  output [15:0] io_deq_bits_31,
  output [1:0]  io_count
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_62;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ram_0 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_1 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_2 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_3 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_4 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_5 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_6 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_7 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_8 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_8_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_8_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_8_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_8_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_8_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_8_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_8_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_9 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_9_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_9_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_9_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_9_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_9_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_9_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_9_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_10 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_10_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_10_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_10_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_10_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_10_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_10_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_10_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_11 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_11_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_11_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_11_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_11_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_11_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_11_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_11_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_12 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_12_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_12_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_12_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_12_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_12_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_12_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_12_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_13 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_13_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_13_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_13_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_13_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_13_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_13_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_13_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_14 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_14_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_14_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_14_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_14_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_14_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_14_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_14_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_15 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_15_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_15_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_15_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_15_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_15_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_15_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_15_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_16 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_16_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_16_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_16_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_16_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_16_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_16_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_16_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_17 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_17_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_17_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_17_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_17_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_17_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_17_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_17_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_18 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_18_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_18_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_18_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_18_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_18_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_18_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_18_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_19 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_19_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_19_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_19_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_19_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_19_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_19_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_19_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_20 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_20_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_20_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_20_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_20_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_20_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_20_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_20_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_21 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_21_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_21_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_21_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_21_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_21_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_21_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_21_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_22 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_22_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_22_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_22_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_22_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_22_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_22_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_22_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_23 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_23_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_23_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_23_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_23_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_23_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_23_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_23_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_24 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_24_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_24_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_24_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_24_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_24_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_24_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_24_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_25 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_25_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_25_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_25_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_25_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_25_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_25_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_25_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_26 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_26_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_26_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_26_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_26_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_26_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_26_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_26_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_27 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_27_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_27_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_27_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_27_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_27_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_27_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_27_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_28 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_28_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_28_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_28_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_28_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_28_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_28_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_28_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_29 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_29_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_29_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_29_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_29_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_29_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_29_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_29_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_30 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_30_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_30_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_30_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_30_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_30_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_30_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_30_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_31 [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_31_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_31_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_31_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_31_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_31_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_31_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_31_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  wrap = enq_ptr_value == 2'h2; // @[Counter.scala 74:24]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  wire  _GEN_45 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_45 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  wrap_1 = deq_ptr_value == 2'h2; // @[Counter.scala 74:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  wire [1:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 312:32]
  wire [1:0] _io_count_T = maybe_full ? 2'h3 : 2'h0; // @[Decoupled.scala 319:10]
  wire [1:0] _io_count_T_3 = 2'h3 + ptr_diff; // @[Decoupled.scala 320:57]
  wire [1:0] _io_count_T_4 = deq_ptr_value > enq_ptr_value ? _io_count_T_3 : ptr_diff; // @[Decoupled.scala 320:10]
  assign ram_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_0_io_deq_bits_MPORT_data = ram_0[ram_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_0_io_deq_bits_MPORT_data = ram_0_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_1[15:0] :
    ram_0[ram_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_0_MPORT_data = io_enq_bits_0;
  assign ram_0_MPORT_addr = enq_ptr_value;
  assign ram_0_MPORT_mask = 1'h1;
  assign ram_0_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_1_io_deq_bits_MPORT_data = ram_1[ram_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_1_io_deq_bits_MPORT_data = ram_1_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_3[15:0] :
    ram_1[ram_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_1_MPORT_data = io_enq_bits_1;
  assign ram_1_MPORT_addr = enq_ptr_value;
  assign ram_1_MPORT_mask = 1'h1;
  assign ram_1_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_2_io_deq_bits_MPORT_data = ram_2[ram_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_2_io_deq_bits_MPORT_data = ram_2_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_5[15:0] :
    ram_2[ram_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_2_MPORT_data = io_enq_bits_2;
  assign ram_2_MPORT_addr = enq_ptr_value;
  assign ram_2_MPORT_mask = 1'h1;
  assign ram_2_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_3_io_deq_bits_MPORT_data = ram_3[ram_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_3_io_deq_bits_MPORT_data = ram_3_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_7[15:0] :
    ram_3[ram_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_3_MPORT_data = io_enq_bits_3;
  assign ram_3_MPORT_addr = enq_ptr_value;
  assign ram_3_MPORT_mask = 1'h1;
  assign ram_3_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_4_io_deq_bits_MPORT_data = ram_4[ram_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_4_io_deq_bits_MPORT_data = ram_4_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_9[15:0] :
    ram_4[ram_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_4_MPORT_data = io_enq_bits_4;
  assign ram_4_MPORT_addr = enq_ptr_value;
  assign ram_4_MPORT_mask = 1'h1;
  assign ram_4_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_5_io_deq_bits_MPORT_data = ram_5[ram_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_5_io_deq_bits_MPORT_data = ram_5_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_11[15:0] :
    ram_5[ram_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_5_MPORT_data = io_enq_bits_5;
  assign ram_5_MPORT_addr = enq_ptr_value;
  assign ram_5_MPORT_mask = 1'h1;
  assign ram_5_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_6_io_deq_bits_MPORT_data = ram_6[ram_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_6_io_deq_bits_MPORT_data = ram_6_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_13[15:0] :
    ram_6[ram_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_6_MPORT_data = io_enq_bits_6;
  assign ram_6_MPORT_addr = enq_ptr_value;
  assign ram_6_MPORT_mask = 1'h1;
  assign ram_6_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_7_io_deq_bits_MPORT_data = ram_7[ram_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_7_io_deq_bits_MPORT_data = ram_7_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_15[15:0] :
    ram_7[ram_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_7_MPORT_data = io_enq_bits_7;
  assign ram_7_MPORT_addr = enq_ptr_value;
  assign ram_7_MPORT_mask = 1'h1;
  assign ram_7_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_8_io_deq_bits_MPORT_en = 1'h1;
  assign ram_8_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_8_io_deq_bits_MPORT_data = ram_8[ram_8_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_8_io_deq_bits_MPORT_data = ram_8_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_17[15:0] :
    ram_8[ram_8_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_8_MPORT_data = io_enq_bits_8;
  assign ram_8_MPORT_addr = enq_ptr_value;
  assign ram_8_MPORT_mask = 1'h1;
  assign ram_8_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_9_io_deq_bits_MPORT_en = 1'h1;
  assign ram_9_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_9_io_deq_bits_MPORT_data = ram_9[ram_9_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_9_io_deq_bits_MPORT_data = ram_9_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_19[15:0] :
    ram_9[ram_9_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_9_MPORT_data = io_enq_bits_9;
  assign ram_9_MPORT_addr = enq_ptr_value;
  assign ram_9_MPORT_mask = 1'h1;
  assign ram_9_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_10_io_deq_bits_MPORT_en = 1'h1;
  assign ram_10_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_10_io_deq_bits_MPORT_data = ram_10[ram_10_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_10_io_deq_bits_MPORT_data = ram_10_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_21[15:0] :
    ram_10[ram_10_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_10_MPORT_data = io_enq_bits_10;
  assign ram_10_MPORT_addr = enq_ptr_value;
  assign ram_10_MPORT_mask = 1'h1;
  assign ram_10_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_11_io_deq_bits_MPORT_en = 1'h1;
  assign ram_11_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_11_io_deq_bits_MPORT_data = ram_11[ram_11_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_11_io_deq_bits_MPORT_data = ram_11_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_23[15:0] :
    ram_11[ram_11_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_11_MPORT_data = io_enq_bits_11;
  assign ram_11_MPORT_addr = enq_ptr_value;
  assign ram_11_MPORT_mask = 1'h1;
  assign ram_11_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_12_io_deq_bits_MPORT_en = 1'h1;
  assign ram_12_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_12_io_deq_bits_MPORT_data = ram_12[ram_12_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_12_io_deq_bits_MPORT_data = ram_12_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_25[15:0] :
    ram_12[ram_12_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_12_MPORT_data = io_enq_bits_12;
  assign ram_12_MPORT_addr = enq_ptr_value;
  assign ram_12_MPORT_mask = 1'h1;
  assign ram_12_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_13_io_deq_bits_MPORT_en = 1'h1;
  assign ram_13_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_13_io_deq_bits_MPORT_data = ram_13[ram_13_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_13_io_deq_bits_MPORT_data = ram_13_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_27[15:0] :
    ram_13[ram_13_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_13_MPORT_data = io_enq_bits_13;
  assign ram_13_MPORT_addr = enq_ptr_value;
  assign ram_13_MPORT_mask = 1'h1;
  assign ram_13_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_14_io_deq_bits_MPORT_en = 1'h1;
  assign ram_14_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_14_io_deq_bits_MPORT_data = ram_14[ram_14_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_14_io_deq_bits_MPORT_data = ram_14_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_29[15:0] :
    ram_14[ram_14_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_14_MPORT_data = io_enq_bits_14;
  assign ram_14_MPORT_addr = enq_ptr_value;
  assign ram_14_MPORT_mask = 1'h1;
  assign ram_14_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_15_io_deq_bits_MPORT_en = 1'h1;
  assign ram_15_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_15_io_deq_bits_MPORT_data = ram_15[ram_15_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_15_io_deq_bits_MPORT_data = ram_15_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_31[15:0] :
    ram_15[ram_15_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_15_MPORT_data = io_enq_bits_15;
  assign ram_15_MPORT_addr = enq_ptr_value;
  assign ram_15_MPORT_mask = 1'h1;
  assign ram_15_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_16_io_deq_bits_MPORT_en = 1'h1;
  assign ram_16_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_16_io_deq_bits_MPORT_data = ram_16[ram_16_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_16_io_deq_bits_MPORT_data = ram_16_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_33[15:0] :
    ram_16[ram_16_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_16_MPORT_data = io_enq_bits_16;
  assign ram_16_MPORT_addr = enq_ptr_value;
  assign ram_16_MPORT_mask = 1'h1;
  assign ram_16_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_17_io_deq_bits_MPORT_en = 1'h1;
  assign ram_17_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_17_io_deq_bits_MPORT_data = ram_17[ram_17_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_17_io_deq_bits_MPORT_data = ram_17_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_35[15:0] :
    ram_17[ram_17_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_17_MPORT_data = io_enq_bits_17;
  assign ram_17_MPORT_addr = enq_ptr_value;
  assign ram_17_MPORT_mask = 1'h1;
  assign ram_17_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_18_io_deq_bits_MPORT_en = 1'h1;
  assign ram_18_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_18_io_deq_bits_MPORT_data = ram_18[ram_18_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_18_io_deq_bits_MPORT_data = ram_18_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_37[15:0] :
    ram_18[ram_18_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_18_MPORT_data = io_enq_bits_18;
  assign ram_18_MPORT_addr = enq_ptr_value;
  assign ram_18_MPORT_mask = 1'h1;
  assign ram_18_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_19_io_deq_bits_MPORT_en = 1'h1;
  assign ram_19_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_19_io_deq_bits_MPORT_data = ram_19[ram_19_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_19_io_deq_bits_MPORT_data = ram_19_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_39[15:0] :
    ram_19[ram_19_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_19_MPORT_data = io_enq_bits_19;
  assign ram_19_MPORT_addr = enq_ptr_value;
  assign ram_19_MPORT_mask = 1'h1;
  assign ram_19_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_20_io_deq_bits_MPORT_en = 1'h1;
  assign ram_20_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_20_io_deq_bits_MPORT_data = ram_20[ram_20_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_20_io_deq_bits_MPORT_data = ram_20_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_41[15:0] :
    ram_20[ram_20_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_20_MPORT_data = io_enq_bits_20;
  assign ram_20_MPORT_addr = enq_ptr_value;
  assign ram_20_MPORT_mask = 1'h1;
  assign ram_20_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_21_io_deq_bits_MPORT_en = 1'h1;
  assign ram_21_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_21_io_deq_bits_MPORT_data = ram_21[ram_21_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_21_io_deq_bits_MPORT_data = ram_21_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_43[15:0] :
    ram_21[ram_21_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_21_MPORT_data = io_enq_bits_21;
  assign ram_21_MPORT_addr = enq_ptr_value;
  assign ram_21_MPORT_mask = 1'h1;
  assign ram_21_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_22_io_deq_bits_MPORT_en = 1'h1;
  assign ram_22_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_22_io_deq_bits_MPORT_data = ram_22[ram_22_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_22_io_deq_bits_MPORT_data = ram_22_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_45[15:0] :
    ram_22[ram_22_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_22_MPORT_data = io_enq_bits_22;
  assign ram_22_MPORT_addr = enq_ptr_value;
  assign ram_22_MPORT_mask = 1'h1;
  assign ram_22_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_23_io_deq_bits_MPORT_en = 1'h1;
  assign ram_23_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_23_io_deq_bits_MPORT_data = ram_23[ram_23_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_23_io_deq_bits_MPORT_data = ram_23_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_47[15:0] :
    ram_23[ram_23_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_23_MPORT_data = io_enq_bits_23;
  assign ram_23_MPORT_addr = enq_ptr_value;
  assign ram_23_MPORT_mask = 1'h1;
  assign ram_23_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_24_io_deq_bits_MPORT_en = 1'h1;
  assign ram_24_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_24_io_deq_bits_MPORT_data = ram_24[ram_24_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_24_io_deq_bits_MPORT_data = ram_24_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_49[15:0] :
    ram_24[ram_24_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_24_MPORT_data = io_enq_bits_24;
  assign ram_24_MPORT_addr = enq_ptr_value;
  assign ram_24_MPORT_mask = 1'h1;
  assign ram_24_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_25_io_deq_bits_MPORT_en = 1'h1;
  assign ram_25_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_25_io_deq_bits_MPORT_data = ram_25[ram_25_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_25_io_deq_bits_MPORT_data = ram_25_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_51[15:0] :
    ram_25[ram_25_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_25_MPORT_data = io_enq_bits_25;
  assign ram_25_MPORT_addr = enq_ptr_value;
  assign ram_25_MPORT_mask = 1'h1;
  assign ram_25_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_26_io_deq_bits_MPORT_en = 1'h1;
  assign ram_26_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_26_io_deq_bits_MPORT_data = ram_26[ram_26_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_26_io_deq_bits_MPORT_data = ram_26_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_53[15:0] :
    ram_26[ram_26_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_26_MPORT_data = io_enq_bits_26;
  assign ram_26_MPORT_addr = enq_ptr_value;
  assign ram_26_MPORT_mask = 1'h1;
  assign ram_26_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_27_io_deq_bits_MPORT_en = 1'h1;
  assign ram_27_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_27_io_deq_bits_MPORT_data = ram_27[ram_27_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_27_io_deq_bits_MPORT_data = ram_27_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_55[15:0] :
    ram_27[ram_27_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_27_MPORT_data = io_enq_bits_27;
  assign ram_27_MPORT_addr = enq_ptr_value;
  assign ram_27_MPORT_mask = 1'h1;
  assign ram_27_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_28_io_deq_bits_MPORT_en = 1'h1;
  assign ram_28_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_28_io_deq_bits_MPORT_data = ram_28[ram_28_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_28_io_deq_bits_MPORT_data = ram_28_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_57[15:0] :
    ram_28[ram_28_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_28_MPORT_data = io_enq_bits_28;
  assign ram_28_MPORT_addr = enq_ptr_value;
  assign ram_28_MPORT_mask = 1'h1;
  assign ram_28_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_29_io_deq_bits_MPORT_en = 1'h1;
  assign ram_29_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_29_io_deq_bits_MPORT_data = ram_29[ram_29_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_29_io_deq_bits_MPORT_data = ram_29_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_59[15:0] :
    ram_29[ram_29_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_29_MPORT_data = io_enq_bits_29;
  assign ram_29_MPORT_addr = enq_ptr_value;
  assign ram_29_MPORT_mask = 1'h1;
  assign ram_29_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_30_io_deq_bits_MPORT_en = 1'h1;
  assign ram_30_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_30_io_deq_bits_MPORT_data = ram_30[ram_30_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_30_io_deq_bits_MPORT_data = ram_30_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_61[15:0] :
    ram_30[ram_30_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_30_MPORT_data = io_enq_bits_30;
  assign ram_30_MPORT_addr = enq_ptr_value;
  assign ram_30_MPORT_mask = 1'h1;
  assign ram_30_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign ram_31_io_deq_bits_MPORT_en = 1'h1;
  assign ram_31_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_31_io_deq_bits_MPORT_data = ram_31[ram_31_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_31_io_deq_bits_MPORT_data = ram_31_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_63[15:0] :
    ram_31[ram_31_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_31_MPORT_data = io_enq_bits_31;
  assign ram_31_MPORT_addr = enq_ptr_value;
  assign ram_31_MPORT_mask = 1'h1;
  assign ram_31_MPORT_en = empty ? _GEN_45 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_0 = empty ? $signed(io_enq_bits_0) : $signed(ram_0_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_1 = empty ? $signed(io_enq_bits_1) : $signed(ram_1_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_2 = empty ? $signed(io_enq_bits_2) : $signed(ram_2_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_3 = empty ? $signed(io_enq_bits_3) : $signed(ram_3_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_4 = empty ? $signed(io_enq_bits_4) : $signed(ram_4_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_5 = empty ? $signed(io_enq_bits_5) : $signed(ram_5_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_6 = empty ? $signed(io_enq_bits_6) : $signed(ram_6_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_7 = empty ? $signed(io_enq_bits_7) : $signed(ram_7_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_8 = empty ? $signed(io_enq_bits_8) : $signed(ram_8_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_9 = empty ? $signed(io_enq_bits_9) : $signed(ram_9_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_10 = empty ? $signed(io_enq_bits_10) : $signed(ram_10_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_11 = empty ? $signed(io_enq_bits_11) : $signed(ram_11_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_12 = empty ? $signed(io_enq_bits_12) : $signed(ram_12_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_13 = empty ? $signed(io_enq_bits_13) : $signed(ram_13_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_14 = empty ? $signed(io_enq_bits_14) : $signed(ram_14_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_15 = empty ? $signed(io_enq_bits_15) : $signed(ram_15_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_16 = empty ? $signed(io_enq_bits_16) : $signed(ram_16_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_17 = empty ? $signed(io_enq_bits_17) : $signed(ram_17_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_18 = empty ? $signed(io_enq_bits_18) : $signed(ram_18_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_19 = empty ? $signed(io_enq_bits_19) : $signed(ram_19_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_20 = empty ? $signed(io_enq_bits_20) : $signed(ram_20_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_21 = empty ? $signed(io_enq_bits_21) : $signed(ram_21_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_22 = empty ? $signed(io_enq_bits_22) : $signed(ram_22_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_23 = empty ? $signed(io_enq_bits_23) : $signed(ram_23_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_24 = empty ? $signed(io_enq_bits_24) : $signed(ram_24_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_25 = empty ? $signed(io_enq_bits_25) : $signed(ram_25_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_26 = empty ? $signed(io_enq_bits_26) : $signed(ram_26_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_27 = empty ? $signed(io_enq_bits_27) : $signed(ram_27_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_28 = empty ? $signed(io_enq_bits_28) : $signed(ram_28_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_29 = empty ? $signed(io_enq_bits_29) : $signed(ram_29_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_30 = empty ? $signed(io_enq_bits_30) : $signed(ram_30_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_31 = empty ? $signed(io_enq_bits_31) : $signed(ram_31_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_count = ptr_match ? _io_count_T : _io_count_T_4; // @[Decoupled.scala 317:20]
  always @(posedge clock) begin
    if (ram_0_MPORT_en & ram_0_MPORT_mask) begin
      ram_0[ram_0_MPORT_addr] <= ram_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_1_MPORT_en & ram_1_MPORT_mask) begin
      ram_1[ram_1_MPORT_addr] <= ram_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_2_MPORT_en & ram_2_MPORT_mask) begin
      ram_2[ram_2_MPORT_addr] <= ram_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_3_MPORT_en & ram_3_MPORT_mask) begin
      ram_3[ram_3_MPORT_addr] <= ram_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_4_MPORT_en & ram_4_MPORT_mask) begin
      ram_4[ram_4_MPORT_addr] <= ram_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_5_MPORT_en & ram_5_MPORT_mask) begin
      ram_5[ram_5_MPORT_addr] <= ram_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_6_MPORT_en & ram_6_MPORT_mask) begin
      ram_6[ram_6_MPORT_addr] <= ram_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_7_MPORT_en & ram_7_MPORT_mask) begin
      ram_7[ram_7_MPORT_addr] <= ram_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_8_MPORT_en & ram_8_MPORT_mask) begin
      ram_8[ram_8_MPORT_addr] <= ram_8_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_9_MPORT_en & ram_9_MPORT_mask) begin
      ram_9[ram_9_MPORT_addr] <= ram_9_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_10_MPORT_en & ram_10_MPORT_mask) begin
      ram_10[ram_10_MPORT_addr] <= ram_10_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_11_MPORT_en & ram_11_MPORT_mask) begin
      ram_11[ram_11_MPORT_addr] <= ram_11_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_12_MPORT_en & ram_12_MPORT_mask) begin
      ram_12[ram_12_MPORT_addr] <= ram_12_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_13_MPORT_en & ram_13_MPORT_mask) begin
      ram_13[ram_13_MPORT_addr] <= ram_13_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_14_MPORT_en & ram_14_MPORT_mask) begin
      ram_14[ram_14_MPORT_addr] <= ram_14_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_15_MPORT_en & ram_15_MPORT_mask) begin
      ram_15[ram_15_MPORT_addr] <= ram_15_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_16_MPORT_en & ram_16_MPORT_mask) begin
      ram_16[ram_16_MPORT_addr] <= ram_16_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_17_MPORT_en & ram_17_MPORT_mask) begin
      ram_17[ram_17_MPORT_addr] <= ram_17_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_18_MPORT_en & ram_18_MPORT_mask) begin
      ram_18[ram_18_MPORT_addr] <= ram_18_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_19_MPORT_en & ram_19_MPORT_mask) begin
      ram_19[ram_19_MPORT_addr] <= ram_19_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_20_MPORT_en & ram_20_MPORT_mask) begin
      ram_20[ram_20_MPORT_addr] <= ram_20_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_21_MPORT_en & ram_21_MPORT_mask) begin
      ram_21[ram_21_MPORT_addr] <= ram_21_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_22_MPORT_en & ram_22_MPORT_mask) begin
      ram_22[ram_22_MPORT_addr] <= ram_22_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_23_MPORT_en & ram_23_MPORT_mask) begin
      ram_23[ram_23_MPORT_addr] <= ram_23_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_24_MPORT_en & ram_24_MPORT_mask) begin
      ram_24[ram_24_MPORT_addr] <= ram_24_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_25_MPORT_en & ram_25_MPORT_mask) begin
      ram_25[ram_25_MPORT_addr] <= ram_25_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_26_MPORT_en & ram_26_MPORT_mask) begin
      ram_26[ram_26_MPORT_addr] <= ram_26_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_27_MPORT_en & ram_27_MPORT_mask) begin
      ram_27[ram_27_MPORT_addr] <= ram_27_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_28_MPORT_en & ram_28_MPORT_mask) begin
      ram_28[ram_28_MPORT_addr] <= ram_28_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_29_MPORT_en & ram_29_MPORT_mask) begin
      ram_29[ram_29_MPORT_addr] <= ram_29_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_30_MPORT_en & ram_30_MPORT_mask) begin
      ram_30[ram_30_MPORT_addr] <= ram_30_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_31_MPORT_en & ram_31_MPORT_mask) begin
      ram_31[ram_31_MPORT_addr] <= ram_31_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      if (wrap) begin // @[Counter.scala 88:20]
        enq_ptr_value <= 2'h0; // @[Counter.scala 88:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      if (wrap_1) begin // @[Counter.scala 88:20]
        deq_ptr_value <= 2'h0; // @[Counter.scala 88:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
  _RAND_17 = {1{`RANDOM}};
  _RAND_19 = {1{`RANDOM}};
  _RAND_21 = {1{`RANDOM}};
  _RAND_23 = {1{`RANDOM}};
  _RAND_25 = {1{`RANDOM}};
  _RAND_27 = {1{`RANDOM}};
  _RAND_29 = {1{`RANDOM}};
  _RAND_31 = {1{`RANDOM}};
  _RAND_33 = {1{`RANDOM}};
  _RAND_35 = {1{`RANDOM}};
  _RAND_37 = {1{`RANDOM}};
  _RAND_39 = {1{`RANDOM}};
  _RAND_41 = {1{`RANDOM}};
  _RAND_43 = {1{`RANDOM}};
  _RAND_45 = {1{`RANDOM}};
  _RAND_47 = {1{`RANDOM}};
  _RAND_49 = {1{`RANDOM}};
  _RAND_51 = {1{`RANDOM}};
  _RAND_53 = {1{`RANDOM}};
  _RAND_55 = {1{`RANDOM}};
  _RAND_57 = {1{`RANDOM}};
  _RAND_59 = {1{`RANDOM}};
  _RAND_61 = {1{`RANDOM}};
  _RAND_63 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_0[initvar] = _RAND_0[15:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_1[initvar] = _RAND_2[15:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_2[initvar] = _RAND_4[15:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_3[initvar] = _RAND_6[15:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_4[initvar] = _RAND_8[15:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_5[initvar] = _RAND_10[15:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_6[initvar] = _RAND_12[15:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_7[initvar] = _RAND_14[15:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_8[initvar] = _RAND_16[15:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_9[initvar] = _RAND_18[15:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_10[initvar] = _RAND_20[15:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_11[initvar] = _RAND_22[15:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_12[initvar] = _RAND_24[15:0];
  _RAND_26 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_13[initvar] = _RAND_26[15:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_14[initvar] = _RAND_28[15:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_15[initvar] = _RAND_30[15:0];
  _RAND_32 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_16[initvar] = _RAND_32[15:0];
  _RAND_34 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_17[initvar] = _RAND_34[15:0];
  _RAND_36 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_18[initvar] = _RAND_36[15:0];
  _RAND_38 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_19[initvar] = _RAND_38[15:0];
  _RAND_40 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_20[initvar] = _RAND_40[15:0];
  _RAND_42 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_21[initvar] = _RAND_42[15:0];
  _RAND_44 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_22[initvar] = _RAND_44[15:0];
  _RAND_46 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_23[initvar] = _RAND_46[15:0];
  _RAND_48 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_24[initvar] = _RAND_48[15:0];
  _RAND_50 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_25[initvar] = _RAND_50[15:0];
  _RAND_52 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_26[initvar] = _RAND_52[15:0];
  _RAND_54 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_27[initvar] = _RAND_54[15:0];
  _RAND_56 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_28[initvar] = _RAND_56[15:0];
  _RAND_58 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_29[initvar] = _RAND_58[15:0];
  _RAND_60 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_30[initvar] = _RAND_60[15:0];
  _RAND_62 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_31[initvar] = _RAND_62[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  enq_ptr_value = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  deq_ptr_value = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  maybe_full = _RAND_66[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualPortMem(
  input         clock,
  input         reset,
  output        io_portA_control_ready,
  input         io_portA_control_valid,
  input         io_portA_control_bits_write,
  input  [11:0] io_portA_control_bits_address,
  output        io_portA_input_ready,
  input         io_portA_input_valid,
  input  [15:0] io_portA_input_bits_0,
  input  [15:0] io_portA_input_bits_1,
  input  [15:0] io_portA_input_bits_2,
  input  [15:0] io_portA_input_bits_3,
  input  [15:0] io_portA_input_bits_4,
  input  [15:0] io_portA_input_bits_5,
  input  [15:0] io_portA_input_bits_6,
  input  [15:0] io_portA_input_bits_7,
  input  [15:0] io_portA_input_bits_8,
  input  [15:0] io_portA_input_bits_9,
  input  [15:0] io_portA_input_bits_10,
  input  [15:0] io_portA_input_bits_11,
  input  [15:0] io_portA_input_bits_12,
  input  [15:0] io_portA_input_bits_13,
  input  [15:0] io_portA_input_bits_14,
  input  [15:0] io_portA_input_bits_15,
  input  [15:0] io_portA_input_bits_16,
  input  [15:0] io_portA_input_bits_17,
  input  [15:0] io_portA_input_bits_18,
  input  [15:0] io_portA_input_bits_19,
  input  [15:0] io_portA_input_bits_20,
  input  [15:0] io_portA_input_bits_21,
  input  [15:0] io_portA_input_bits_22,
  input  [15:0] io_portA_input_bits_23,
  input  [15:0] io_portA_input_bits_24,
  input  [15:0] io_portA_input_bits_25,
  input  [15:0] io_portA_input_bits_26,
  input  [15:0] io_portA_input_bits_27,
  input  [15:0] io_portA_input_bits_28,
  input  [15:0] io_portA_input_bits_29,
  input  [15:0] io_portA_input_bits_30,
  input  [15:0] io_portA_input_bits_31,
  input         io_portA_output_ready,
  output        io_portA_output_valid,
  output [15:0] io_portA_output_bits_0,
  output [15:0] io_portA_output_bits_1,
  output [15:0] io_portA_output_bits_2,
  output [15:0] io_portA_output_bits_3,
  output [15:0] io_portA_output_bits_4,
  output [15:0] io_portA_output_bits_5,
  output [15:0] io_portA_output_bits_6,
  output [15:0] io_portA_output_bits_7,
  output [15:0] io_portA_output_bits_8,
  output [15:0] io_portA_output_bits_9,
  output [15:0] io_portA_output_bits_10,
  output [15:0] io_portA_output_bits_11,
  output [15:0] io_portA_output_bits_12,
  output [15:0] io_portA_output_bits_13,
  output [15:0] io_portA_output_bits_14,
  output [15:0] io_portA_output_bits_15,
  output [15:0] io_portA_output_bits_16,
  output [15:0] io_portA_output_bits_17,
  output [15:0] io_portA_output_bits_18,
  output [15:0] io_portA_output_bits_19,
  output [15:0] io_portA_output_bits_20,
  output [15:0] io_portA_output_bits_21,
  output [15:0] io_portA_output_bits_22,
  output [15:0] io_portA_output_bits_23,
  output [15:0] io_portA_output_bits_24,
  output [15:0] io_portA_output_bits_25,
  output [15:0] io_portA_output_bits_26,
  output [15:0] io_portA_output_bits_27,
  output [15:0] io_portA_output_bits_28,
  output [15:0] io_portA_output_bits_29,
  output [15:0] io_portA_output_bits_30,
  output [15:0] io_portA_output_bits_31,
  output        io_portB_control_ready,
  input         io_portB_control_valid,
  input  [11:0] io_portB_control_bits_address,
  input         io_portB_output_ready,
  output        io_portB_output_valid,
  output [15:0] io_portB_output_bits_0,
  output [15:0] io_portB_output_bits_1,
  output [15:0] io_portB_output_bits_2,
  output [15:0] io_portB_output_bits_3,
  output [15:0] io_portB_output_bits_4,
  output [15:0] io_portB_output_bits_5,
  output [15:0] io_portB_output_bits_6,
  output [15:0] io_portB_output_bits_7,
  output [15:0] io_portB_output_bits_8,
  output [15:0] io_portB_output_bits_9,
  output [15:0] io_portB_output_bits_10,
  output [15:0] io_portB_output_bits_11,
  output [15:0] io_portB_output_bits_12,
  output [15:0] io_portB_output_bits_13,
  output [15:0] io_portB_output_bits_14,
  output [15:0] io_portB_output_bits_15,
  output [15:0] io_portB_output_bits_16,
  output [15:0] io_portB_output_bits_17,
  output [15:0] io_portB_output_bits_18,
  output [15:0] io_portB_output_bits_19,
  output [15:0] io_portB_output_bits_20,
  output [15:0] io_portB_output_bits_21,
  output [15:0] io_portB_output_bits_22,
  output [15:0] io_portB_output_bits_23,
  output [15:0] io_portB_output_bits_24,
  output [15:0] io_portB_output_bits_25,
  output [15:0] io_portB_output_bits_26,
  output [15:0] io_portB_output_bits_27,
  output [15:0] io_portB_output_bits_28,
  output [15:0] io_portB_output_bits_29,
  output [15:0] io_portB_output_bits_30,
  output [15:0] io_portB_output_bits_31,
  input         io_tracepoint,
  input  [31:0] io_programCounter
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  mem_clock; // @[DualPortMem.scala 33:19]
  wire  mem_reset; // @[DualPortMem.scala 33:19]
  wire [11:0] mem_io_portA_address; // @[DualPortMem.scala 33:19]
  wire  mem_io_portA_read_enable; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_0; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_1; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_2; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_3; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_4; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_5; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_6; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_7; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_8; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_9; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_10; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_11; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_12; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_13; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_14; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_15; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_16; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_17; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_18; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_19; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_20; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_21; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_22; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_23; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_24; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_25; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_26; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_27; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_28; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_29; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_30; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_31; // @[DualPortMem.scala 33:19]
  wire  mem_io_portA_write_enable; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_0; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_1; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_2; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_3; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_4; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_5; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_6; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_7; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_8; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_9; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_10; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_11; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_12; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_13; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_14; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_15; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_16; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_17; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_18; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_19; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_20; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_21; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_22; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_23; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_24; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_25; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_26; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_27; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_28; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_29; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_30; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_31; // @[DualPortMem.scala 33:19]
  wire [11:0] mem_io_portB_address; // @[DualPortMem.scala 33:19]
  wire  mem_io_portB_read_enable; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_0; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_1; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_2; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_3; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_4; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_5; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_6; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_7; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_8; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_9; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_10; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_11; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_12; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_13; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_14; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_15; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_16; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_17; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_18; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_19; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_20; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_21; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_22; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_23; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_24; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_25; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_26; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_27; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_28; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_29; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_30; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_31; // @[DualPortMem.scala 33:19]
  wire  output__clock; // @[DualPortMem.scala 48:24]
  wire  output__reset; // @[DualPortMem.scala 48:24]
  wire  output__io_enq_ready; // @[DualPortMem.scala 48:24]
  wire  output__io_enq_valid; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_0; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_1; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_2; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_3; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_4; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_5; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_6; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_7; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_8; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_9; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_10; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_11; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_12; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_13; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_14; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_15; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_16; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_17; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_18; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_19; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_20; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_21; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_22; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_23; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_24; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_25; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_26; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_27; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_28; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_29; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_30; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_31; // @[DualPortMem.scala 48:24]
  wire  output__io_deq_ready; // @[DualPortMem.scala 48:24]
  wire  output__io_deq_valid; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_0; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_1; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_2; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_3; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_4; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_5; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_6; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_7; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_8; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_9; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_10; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_11; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_12; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_13; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_14; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_15; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_16; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_17; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_18; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_19; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_20; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_21; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_22; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_23; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_24; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_25; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_26; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_27; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_28; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_29; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_30; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_31; // @[DualPortMem.scala 48:24]
  wire [1:0] output__io_count; // @[DualPortMem.scala 48:24]
  wire  output_1_clock; // @[DualPortMem.scala 48:24]
  wire  output_1_reset; // @[DualPortMem.scala 48:24]
  wire  output_1_io_enq_ready; // @[DualPortMem.scala 48:24]
  wire  output_1_io_enq_valid; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_0; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_1; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_2; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_3; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_4; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_5; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_6; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_7; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_8; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_9; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_10; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_11; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_12; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_13; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_14; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_15; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_16; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_17; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_18; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_19; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_20; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_21; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_22; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_23; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_24; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_25; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_26; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_27; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_28; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_29; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_30; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_31; // @[DualPortMem.scala 48:24]
  wire  output_1_io_deq_ready; // @[DualPortMem.scala 48:24]
  wire  output_1_io_deq_valid; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_0; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_1; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_2; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_3; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_4; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_5; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_6; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_7; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_8; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_9; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_10; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_11; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_12; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_13; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_14; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_15; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_16; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_17; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_18; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_19; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_20; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_21; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_22; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_23; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_24; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_25; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_26; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_27; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_28; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_29; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_30; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_31; // @[DualPortMem.scala 48:24]
  wire [1:0] output_1_io_count; // @[DualPortMem.scala 48:24]
  wire  outputReady = output__io_count < 2'h2; // @[DualPortMem.scala 55:39]
  reg  output_io_enq_valid_sr_0; // @[ShiftRegister.scala 10:22]
  wire  outputReady_1 = output_1_io_count < 2'h2; // @[DualPortMem.scala 55:39]
  reg  output_io_enq_valid_sr_1_0; // @[ShiftRegister.scala 10:22]
  InnerDualPortMem mem ( // @[DualPortMem.scala 33:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_portA_address(mem_io_portA_address),
    .io_portA_read_enable(mem_io_portA_read_enable),
    .io_portA_read_data_0(mem_io_portA_read_data_0),
    .io_portA_read_data_1(mem_io_portA_read_data_1),
    .io_portA_read_data_2(mem_io_portA_read_data_2),
    .io_portA_read_data_3(mem_io_portA_read_data_3),
    .io_portA_read_data_4(mem_io_portA_read_data_4),
    .io_portA_read_data_5(mem_io_portA_read_data_5),
    .io_portA_read_data_6(mem_io_portA_read_data_6),
    .io_portA_read_data_7(mem_io_portA_read_data_7),
    .io_portA_read_data_8(mem_io_portA_read_data_8),
    .io_portA_read_data_9(mem_io_portA_read_data_9),
    .io_portA_read_data_10(mem_io_portA_read_data_10),
    .io_portA_read_data_11(mem_io_portA_read_data_11),
    .io_portA_read_data_12(mem_io_portA_read_data_12),
    .io_portA_read_data_13(mem_io_portA_read_data_13),
    .io_portA_read_data_14(mem_io_portA_read_data_14),
    .io_portA_read_data_15(mem_io_portA_read_data_15),
    .io_portA_read_data_16(mem_io_portA_read_data_16),
    .io_portA_read_data_17(mem_io_portA_read_data_17),
    .io_portA_read_data_18(mem_io_portA_read_data_18),
    .io_portA_read_data_19(mem_io_portA_read_data_19),
    .io_portA_read_data_20(mem_io_portA_read_data_20),
    .io_portA_read_data_21(mem_io_portA_read_data_21),
    .io_portA_read_data_22(mem_io_portA_read_data_22),
    .io_portA_read_data_23(mem_io_portA_read_data_23),
    .io_portA_read_data_24(mem_io_portA_read_data_24),
    .io_portA_read_data_25(mem_io_portA_read_data_25),
    .io_portA_read_data_26(mem_io_portA_read_data_26),
    .io_portA_read_data_27(mem_io_portA_read_data_27),
    .io_portA_read_data_28(mem_io_portA_read_data_28),
    .io_portA_read_data_29(mem_io_portA_read_data_29),
    .io_portA_read_data_30(mem_io_portA_read_data_30),
    .io_portA_read_data_31(mem_io_portA_read_data_31),
    .io_portA_write_enable(mem_io_portA_write_enable),
    .io_portA_write_data_0(mem_io_portA_write_data_0),
    .io_portA_write_data_1(mem_io_portA_write_data_1),
    .io_portA_write_data_2(mem_io_portA_write_data_2),
    .io_portA_write_data_3(mem_io_portA_write_data_3),
    .io_portA_write_data_4(mem_io_portA_write_data_4),
    .io_portA_write_data_5(mem_io_portA_write_data_5),
    .io_portA_write_data_6(mem_io_portA_write_data_6),
    .io_portA_write_data_7(mem_io_portA_write_data_7),
    .io_portA_write_data_8(mem_io_portA_write_data_8),
    .io_portA_write_data_9(mem_io_portA_write_data_9),
    .io_portA_write_data_10(mem_io_portA_write_data_10),
    .io_portA_write_data_11(mem_io_portA_write_data_11),
    .io_portA_write_data_12(mem_io_portA_write_data_12),
    .io_portA_write_data_13(mem_io_portA_write_data_13),
    .io_portA_write_data_14(mem_io_portA_write_data_14),
    .io_portA_write_data_15(mem_io_portA_write_data_15),
    .io_portA_write_data_16(mem_io_portA_write_data_16),
    .io_portA_write_data_17(mem_io_portA_write_data_17),
    .io_portA_write_data_18(mem_io_portA_write_data_18),
    .io_portA_write_data_19(mem_io_portA_write_data_19),
    .io_portA_write_data_20(mem_io_portA_write_data_20),
    .io_portA_write_data_21(mem_io_portA_write_data_21),
    .io_portA_write_data_22(mem_io_portA_write_data_22),
    .io_portA_write_data_23(mem_io_portA_write_data_23),
    .io_portA_write_data_24(mem_io_portA_write_data_24),
    .io_portA_write_data_25(mem_io_portA_write_data_25),
    .io_portA_write_data_26(mem_io_portA_write_data_26),
    .io_portA_write_data_27(mem_io_portA_write_data_27),
    .io_portA_write_data_28(mem_io_portA_write_data_28),
    .io_portA_write_data_29(mem_io_portA_write_data_29),
    .io_portA_write_data_30(mem_io_portA_write_data_30),
    .io_portA_write_data_31(mem_io_portA_write_data_31),
    .io_portB_address(mem_io_portB_address),
    .io_portB_read_enable(mem_io_portB_read_enable),
    .io_portB_read_data_0(mem_io_portB_read_data_0),
    .io_portB_read_data_1(mem_io_portB_read_data_1),
    .io_portB_read_data_2(mem_io_portB_read_data_2),
    .io_portB_read_data_3(mem_io_portB_read_data_3),
    .io_portB_read_data_4(mem_io_portB_read_data_4),
    .io_portB_read_data_5(mem_io_portB_read_data_5),
    .io_portB_read_data_6(mem_io_portB_read_data_6),
    .io_portB_read_data_7(mem_io_portB_read_data_7),
    .io_portB_read_data_8(mem_io_portB_read_data_8),
    .io_portB_read_data_9(mem_io_portB_read_data_9),
    .io_portB_read_data_10(mem_io_portB_read_data_10),
    .io_portB_read_data_11(mem_io_portB_read_data_11),
    .io_portB_read_data_12(mem_io_portB_read_data_12),
    .io_portB_read_data_13(mem_io_portB_read_data_13),
    .io_portB_read_data_14(mem_io_portB_read_data_14),
    .io_portB_read_data_15(mem_io_portB_read_data_15),
    .io_portB_read_data_16(mem_io_portB_read_data_16),
    .io_portB_read_data_17(mem_io_portB_read_data_17),
    .io_portB_read_data_18(mem_io_portB_read_data_18),
    .io_portB_read_data_19(mem_io_portB_read_data_19),
    .io_portB_read_data_20(mem_io_portB_read_data_20),
    .io_portB_read_data_21(mem_io_portB_read_data_21),
    .io_portB_read_data_22(mem_io_portB_read_data_22),
    .io_portB_read_data_23(mem_io_portB_read_data_23),
    .io_portB_read_data_24(mem_io_portB_read_data_24),
    .io_portB_read_data_25(mem_io_portB_read_data_25),
    .io_portB_read_data_26(mem_io_portB_read_data_26),
    .io_portB_read_data_27(mem_io_portB_read_data_27),
    .io_portB_read_data_28(mem_io_portB_read_data_28),
    .io_portB_read_data_29(mem_io_portB_read_data_29),
    .io_portB_read_data_30(mem_io_portB_read_data_30),
    .io_portB_read_data_31(mem_io_portB_read_data_31)
  );
  Queue_10 output_ ( // @[DualPortMem.scala 48:24]
    .clock(output__clock),
    .reset(output__reset),
    .io_enq_ready(output__io_enq_ready),
    .io_enq_valid(output__io_enq_valid),
    .io_enq_bits_0(output__io_enq_bits_0),
    .io_enq_bits_1(output__io_enq_bits_1),
    .io_enq_bits_2(output__io_enq_bits_2),
    .io_enq_bits_3(output__io_enq_bits_3),
    .io_enq_bits_4(output__io_enq_bits_4),
    .io_enq_bits_5(output__io_enq_bits_5),
    .io_enq_bits_6(output__io_enq_bits_6),
    .io_enq_bits_7(output__io_enq_bits_7),
    .io_enq_bits_8(output__io_enq_bits_8),
    .io_enq_bits_9(output__io_enq_bits_9),
    .io_enq_bits_10(output__io_enq_bits_10),
    .io_enq_bits_11(output__io_enq_bits_11),
    .io_enq_bits_12(output__io_enq_bits_12),
    .io_enq_bits_13(output__io_enq_bits_13),
    .io_enq_bits_14(output__io_enq_bits_14),
    .io_enq_bits_15(output__io_enq_bits_15),
    .io_enq_bits_16(output__io_enq_bits_16),
    .io_enq_bits_17(output__io_enq_bits_17),
    .io_enq_bits_18(output__io_enq_bits_18),
    .io_enq_bits_19(output__io_enq_bits_19),
    .io_enq_bits_20(output__io_enq_bits_20),
    .io_enq_bits_21(output__io_enq_bits_21),
    .io_enq_bits_22(output__io_enq_bits_22),
    .io_enq_bits_23(output__io_enq_bits_23),
    .io_enq_bits_24(output__io_enq_bits_24),
    .io_enq_bits_25(output__io_enq_bits_25),
    .io_enq_bits_26(output__io_enq_bits_26),
    .io_enq_bits_27(output__io_enq_bits_27),
    .io_enq_bits_28(output__io_enq_bits_28),
    .io_enq_bits_29(output__io_enq_bits_29),
    .io_enq_bits_30(output__io_enq_bits_30),
    .io_enq_bits_31(output__io_enq_bits_31),
    .io_deq_ready(output__io_deq_ready),
    .io_deq_valid(output__io_deq_valid),
    .io_deq_bits_0(output__io_deq_bits_0),
    .io_deq_bits_1(output__io_deq_bits_1),
    .io_deq_bits_2(output__io_deq_bits_2),
    .io_deq_bits_3(output__io_deq_bits_3),
    .io_deq_bits_4(output__io_deq_bits_4),
    .io_deq_bits_5(output__io_deq_bits_5),
    .io_deq_bits_6(output__io_deq_bits_6),
    .io_deq_bits_7(output__io_deq_bits_7),
    .io_deq_bits_8(output__io_deq_bits_8),
    .io_deq_bits_9(output__io_deq_bits_9),
    .io_deq_bits_10(output__io_deq_bits_10),
    .io_deq_bits_11(output__io_deq_bits_11),
    .io_deq_bits_12(output__io_deq_bits_12),
    .io_deq_bits_13(output__io_deq_bits_13),
    .io_deq_bits_14(output__io_deq_bits_14),
    .io_deq_bits_15(output__io_deq_bits_15),
    .io_deq_bits_16(output__io_deq_bits_16),
    .io_deq_bits_17(output__io_deq_bits_17),
    .io_deq_bits_18(output__io_deq_bits_18),
    .io_deq_bits_19(output__io_deq_bits_19),
    .io_deq_bits_20(output__io_deq_bits_20),
    .io_deq_bits_21(output__io_deq_bits_21),
    .io_deq_bits_22(output__io_deq_bits_22),
    .io_deq_bits_23(output__io_deq_bits_23),
    .io_deq_bits_24(output__io_deq_bits_24),
    .io_deq_bits_25(output__io_deq_bits_25),
    .io_deq_bits_26(output__io_deq_bits_26),
    .io_deq_bits_27(output__io_deq_bits_27),
    .io_deq_bits_28(output__io_deq_bits_28),
    .io_deq_bits_29(output__io_deq_bits_29),
    .io_deq_bits_30(output__io_deq_bits_30),
    .io_deq_bits_31(output__io_deq_bits_31),
    .io_count(output__io_count)
  );
  Queue_10 output_1 ( // @[DualPortMem.scala 48:24]
    .clock(output_1_clock),
    .reset(output_1_reset),
    .io_enq_ready(output_1_io_enq_ready),
    .io_enq_valid(output_1_io_enq_valid),
    .io_enq_bits_0(output_1_io_enq_bits_0),
    .io_enq_bits_1(output_1_io_enq_bits_1),
    .io_enq_bits_2(output_1_io_enq_bits_2),
    .io_enq_bits_3(output_1_io_enq_bits_3),
    .io_enq_bits_4(output_1_io_enq_bits_4),
    .io_enq_bits_5(output_1_io_enq_bits_5),
    .io_enq_bits_6(output_1_io_enq_bits_6),
    .io_enq_bits_7(output_1_io_enq_bits_7),
    .io_enq_bits_8(output_1_io_enq_bits_8),
    .io_enq_bits_9(output_1_io_enq_bits_9),
    .io_enq_bits_10(output_1_io_enq_bits_10),
    .io_enq_bits_11(output_1_io_enq_bits_11),
    .io_enq_bits_12(output_1_io_enq_bits_12),
    .io_enq_bits_13(output_1_io_enq_bits_13),
    .io_enq_bits_14(output_1_io_enq_bits_14),
    .io_enq_bits_15(output_1_io_enq_bits_15),
    .io_enq_bits_16(output_1_io_enq_bits_16),
    .io_enq_bits_17(output_1_io_enq_bits_17),
    .io_enq_bits_18(output_1_io_enq_bits_18),
    .io_enq_bits_19(output_1_io_enq_bits_19),
    .io_enq_bits_20(output_1_io_enq_bits_20),
    .io_enq_bits_21(output_1_io_enq_bits_21),
    .io_enq_bits_22(output_1_io_enq_bits_22),
    .io_enq_bits_23(output_1_io_enq_bits_23),
    .io_enq_bits_24(output_1_io_enq_bits_24),
    .io_enq_bits_25(output_1_io_enq_bits_25),
    .io_enq_bits_26(output_1_io_enq_bits_26),
    .io_enq_bits_27(output_1_io_enq_bits_27),
    .io_enq_bits_28(output_1_io_enq_bits_28),
    .io_enq_bits_29(output_1_io_enq_bits_29),
    .io_enq_bits_30(output_1_io_enq_bits_30),
    .io_enq_bits_31(output_1_io_enq_bits_31),
    .io_deq_ready(output_1_io_deq_ready),
    .io_deq_valid(output_1_io_deq_valid),
    .io_deq_bits_0(output_1_io_deq_bits_0),
    .io_deq_bits_1(output_1_io_deq_bits_1),
    .io_deq_bits_2(output_1_io_deq_bits_2),
    .io_deq_bits_3(output_1_io_deq_bits_3),
    .io_deq_bits_4(output_1_io_deq_bits_4),
    .io_deq_bits_5(output_1_io_deq_bits_5),
    .io_deq_bits_6(output_1_io_deq_bits_6),
    .io_deq_bits_7(output_1_io_deq_bits_7),
    .io_deq_bits_8(output_1_io_deq_bits_8),
    .io_deq_bits_9(output_1_io_deq_bits_9),
    .io_deq_bits_10(output_1_io_deq_bits_10),
    .io_deq_bits_11(output_1_io_deq_bits_11),
    .io_deq_bits_12(output_1_io_deq_bits_12),
    .io_deq_bits_13(output_1_io_deq_bits_13),
    .io_deq_bits_14(output_1_io_deq_bits_14),
    .io_deq_bits_15(output_1_io_deq_bits_15),
    .io_deq_bits_16(output_1_io_deq_bits_16),
    .io_deq_bits_17(output_1_io_deq_bits_17),
    .io_deq_bits_18(output_1_io_deq_bits_18),
    .io_deq_bits_19(output_1_io_deq_bits_19),
    .io_deq_bits_20(output_1_io_deq_bits_20),
    .io_deq_bits_21(output_1_io_deq_bits_21),
    .io_deq_bits_22(output_1_io_deq_bits_22),
    .io_deq_bits_23(output_1_io_deq_bits_23),
    .io_deq_bits_24(output_1_io_deq_bits_24),
    .io_deq_bits_25(output_1_io_deq_bits_25),
    .io_deq_bits_26(output_1_io_deq_bits_26),
    .io_deq_bits_27(output_1_io_deq_bits_27),
    .io_deq_bits_28(output_1_io_deq_bits_28),
    .io_deq_bits_29(output_1_io_deq_bits_29),
    .io_deq_bits_30(output_1_io_deq_bits_30),
    .io_deq_bits_31(output_1_io_deq_bits_31),
    .io_count(output_1_io_count)
  );
  assign io_portA_control_ready = io_portA_control_bits_write ? io_portA_input_valid : outputReady; // @[DualPortMem.scala 59:30 60:21 64:21]
  assign io_portA_input_ready = io_portA_control_valid & io_portA_control_bits_write; // @[DualPortMem.scala 75:34]
  assign io_portA_output_valid = output__io_deq_valid; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_0 = output__io_deq_bits_0; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_1 = output__io_deq_bits_1; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_2 = output__io_deq_bits_2; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_3 = output__io_deq_bits_3; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_4 = output__io_deq_bits_4; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_5 = output__io_deq_bits_5; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_6 = output__io_deq_bits_6; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_7 = output__io_deq_bits_7; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_8 = output__io_deq_bits_8; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_9 = output__io_deq_bits_9; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_10 = output__io_deq_bits_10; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_11 = output__io_deq_bits_11; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_12 = output__io_deq_bits_12; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_13 = output__io_deq_bits_13; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_14 = output__io_deq_bits_14; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_15 = output__io_deq_bits_15; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_16 = output__io_deq_bits_16; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_17 = output__io_deq_bits_17; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_18 = output__io_deq_bits_18; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_19 = output__io_deq_bits_19; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_20 = output__io_deq_bits_20; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_21 = output__io_deq_bits_21; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_22 = output__io_deq_bits_22; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_23 = output__io_deq_bits_23; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_24 = output__io_deq_bits_24; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_25 = output__io_deq_bits_25; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_26 = output__io_deq_bits_26; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_27 = output__io_deq_bits_27; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_28 = output__io_deq_bits_28; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_29 = output__io_deq_bits_29; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_30 = output__io_deq_bits_30; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_31 = output__io_deq_bits_31; // @[DualPortMem.scala 72:17]
  assign io_portB_control_ready = output_1_io_count < 2'h2; // @[DualPortMem.scala 55:39]
  assign io_portB_output_valid = output_1_io_deq_valid; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_0 = output_1_io_deq_bits_0; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_1 = output_1_io_deq_bits_1; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_2 = output_1_io_deq_bits_2; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_3 = output_1_io_deq_bits_3; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_4 = output_1_io_deq_bits_4; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_5 = output_1_io_deq_bits_5; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_6 = output_1_io_deq_bits_6; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_7 = output_1_io_deq_bits_7; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_8 = output_1_io_deq_bits_8; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_9 = output_1_io_deq_bits_9; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_10 = output_1_io_deq_bits_10; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_11 = output_1_io_deq_bits_11; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_12 = output_1_io_deq_bits_12; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_13 = output_1_io_deq_bits_13; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_14 = output_1_io_deq_bits_14; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_15 = output_1_io_deq_bits_15; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_16 = output_1_io_deq_bits_16; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_17 = output_1_io_deq_bits_17; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_18 = output_1_io_deq_bits_18; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_19 = output_1_io_deq_bits_19; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_20 = output_1_io_deq_bits_20; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_21 = output_1_io_deq_bits_21; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_22 = output_1_io_deq_bits_22; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_23 = output_1_io_deq_bits_23; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_24 = output_1_io_deq_bits_24; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_25 = output_1_io_deq_bits_25; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_26 = output_1_io_deq_bits_26; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_27 = output_1_io_deq_bits_27; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_28 = output_1_io_deq_bits_28; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_29 = output_1_io_deq_bits_29; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_30 = output_1_io_deq_bits_30; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_31 = output_1_io_deq_bits_31; // @[DualPortMem.scala 72:17]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_portA_address = io_portA_control_bits_address; // @[DualPortMem.scala 57:19]
  assign mem_io_portA_read_enable = io_portA_control_bits_write ? 1'h0 : io_portA_control_valid & outputReady; // @[DualPortMem.scala 59:30 62:25 66:25]
  assign mem_io_portA_write_enable = io_portA_control_bits_write & (io_portA_control_valid & io_portA_input_valid); // @[DualPortMem.scala 59:30 61:26 65:26]
  assign mem_io_portA_write_data_0 = io_portA_input_bits_0; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_1 = io_portA_input_bits_1; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_2 = io_portA_input_bits_2; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_3 = io_portA_input_bits_3; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_4 = io_portA_input_bits_4; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_5 = io_portA_input_bits_5; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_6 = io_portA_input_bits_6; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_7 = io_portA_input_bits_7; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_8 = io_portA_input_bits_8; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_9 = io_portA_input_bits_9; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_10 = io_portA_input_bits_10; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_11 = io_portA_input_bits_11; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_12 = io_portA_input_bits_12; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_13 = io_portA_input_bits_13; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_14 = io_portA_input_bits_14; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_15 = io_portA_input_bits_15; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_16 = io_portA_input_bits_16; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_17 = io_portA_input_bits_17; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_18 = io_portA_input_bits_18; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_19 = io_portA_input_bits_19; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_20 = io_portA_input_bits_20; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_21 = io_portA_input_bits_21; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_22 = io_portA_input_bits_22; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_23 = io_portA_input_bits_23; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_24 = io_portA_input_bits_24; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_25 = io_portA_input_bits_25; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_26 = io_portA_input_bits_26; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_27 = io_portA_input_bits_27; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_28 = io_portA_input_bits_28; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_29 = io_portA_input_bits_29; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_30 = io_portA_input_bits_30; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_31 = io_portA_input_bits_31; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_address = io_portB_control_bits_address; // @[DualPortMem.scala 57:19]
  assign mem_io_portB_read_enable = io_portB_control_valid & outputReady_1; // @[DualPortMem.scala 66:42]
  assign output__clock = clock;
  assign output__reset = reset;
  assign output__io_enq_valid = output_io_enq_valid_sr_0; // @[DualPortMem.scala 70:25]
  assign output__io_enq_bits_0 = mem_io_portA_read_data_0; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_1 = mem_io_portA_read_data_1; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_2 = mem_io_portA_read_data_2; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_3 = mem_io_portA_read_data_3; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_4 = mem_io_portA_read_data_4; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_5 = mem_io_portA_read_data_5; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_6 = mem_io_portA_read_data_6; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_7 = mem_io_portA_read_data_7; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_8 = mem_io_portA_read_data_8; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_9 = mem_io_portA_read_data_9; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_10 = mem_io_portA_read_data_10; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_11 = mem_io_portA_read_data_11; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_12 = mem_io_portA_read_data_12; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_13 = mem_io_portA_read_data_13; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_14 = mem_io_portA_read_data_14; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_15 = mem_io_portA_read_data_15; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_16 = mem_io_portA_read_data_16; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_17 = mem_io_portA_read_data_17; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_18 = mem_io_portA_read_data_18; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_19 = mem_io_portA_read_data_19; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_20 = mem_io_portA_read_data_20; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_21 = mem_io_portA_read_data_21; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_22 = mem_io_portA_read_data_22; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_23 = mem_io_portA_read_data_23; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_24 = mem_io_portA_read_data_24; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_25 = mem_io_portA_read_data_25; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_26 = mem_io_portA_read_data_26; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_27 = mem_io_portA_read_data_27; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_28 = mem_io_portA_read_data_28; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_29 = mem_io_portA_read_data_29; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_30 = mem_io_portA_read_data_30; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_31 = mem_io_portA_read_data_31; // @[DualPortMem.scala 69:24]
  assign output__io_deq_ready = io_portA_output_ready; // @[DualPortMem.scala 72:17]
  assign output_1_clock = clock;
  assign output_1_reset = reset;
  assign output_1_io_enq_valid = output_io_enq_valid_sr_1_0; // @[DualPortMem.scala 70:25]
  assign output_1_io_enq_bits_0 = mem_io_portB_read_data_0; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_1 = mem_io_portB_read_data_1; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_2 = mem_io_portB_read_data_2; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_3 = mem_io_portB_read_data_3; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_4 = mem_io_portB_read_data_4; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_5 = mem_io_portB_read_data_5; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_6 = mem_io_portB_read_data_6; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_7 = mem_io_portB_read_data_7; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_8 = mem_io_portB_read_data_8; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_9 = mem_io_portB_read_data_9; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_10 = mem_io_portB_read_data_10; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_11 = mem_io_portB_read_data_11; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_12 = mem_io_portB_read_data_12; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_13 = mem_io_portB_read_data_13; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_14 = mem_io_portB_read_data_14; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_15 = mem_io_portB_read_data_15; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_16 = mem_io_portB_read_data_16; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_17 = mem_io_portB_read_data_17; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_18 = mem_io_portB_read_data_18; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_19 = mem_io_portB_read_data_19; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_20 = mem_io_portB_read_data_20; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_21 = mem_io_portB_read_data_21; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_22 = mem_io_portB_read_data_22; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_23 = mem_io_portB_read_data_23; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_24 = mem_io_portB_read_data_24; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_25 = mem_io_portB_read_data_25; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_26 = mem_io_portB_read_data_26; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_27 = mem_io_portB_read_data_27; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_28 = mem_io_portB_read_data_28; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_29 = mem_io_portB_read_data_29; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_30 = mem_io_portB_read_data_30; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_31 = mem_io_portB_read_data_31; // @[DualPortMem.scala 69:24]
  assign output_1_io_deq_ready = io_portB_output_ready; // @[DualPortMem.scala 72:17]
  always @(posedge clock) begin
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_0 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_0 <= mem_io_portA_read_enable; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_1_0 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_1_0 <= mem_io_portB_read_enable; // @[ShiftRegister.scala 25:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  output_io_enq_valid_sr_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  output_io_enq_valid_sr_1_0 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module VecAdder(
  output        io_left_ready,
  input         io_left_valid,
  input  [15:0] io_left_bits_0,
  input  [15:0] io_left_bits_1,
  input  [15:0] io_left_bits_2,
  input  [15:0] io_left_bits_3,
  input  [15:0] io_left_bits_4,
  input  [15:0] io_left_bits_5,
  input  [15:0] io_left_bits_6,
  input  [15:0] io_left_bits_7,
  input  [15:0] io_left_bits_8,
  input  [15:0] io_left_bits_9,
  input  [15:0] io_left_bits_10,
  input  [15:0] io_left_bits_11,
  input  [15:0] io_left_bits_12,
  input  [15:0] io_left_bits_13,
  input  [15:0] io_left_bits_14,
  input  [15:0] io_left_bits_15,
  input  [15:0] io_left_bits_16,
  input  [15:0] io_left_bits_17,
  input  [15:0] io_left_bits_18,
  input  [15:0] io_left_bits_19,
  input  [15:0] io_left_bits_20,
  input  [15:0] io_left_bits_21,
  input  [15:0] io_left_bits_22,
  input  [15:0] io_left_bits_23,
  input  [15:0] io_left_bits_24,
  input  [15:0] io_left_bits_25,
  input  [15:0] io_left_bits_26,
  input  [15:0] io_left_bits_27,
  input  [15:0] io_left_bits_28,
  input  [15:0] io_left_bits_29,
  input  [15:0] io_left_bits_30,
  input  [15:0] io_left_bits_31,
  output        io_right_ready,
  input         io_right_valid,
  input  [15:0] io_right_bits_0,
  input  [15:0] io_right_bits_1,
  input  [15:0] io_right_bits_2,
  input  [15:0] io_right_bits_3,
  input  [15:0] io_right_bits_4,
  input  [15:0] io_right_bits_5,
  input  [15:0] io_right_bits_6,
  input  [15:0] io_right_bits_7,
  input  [15:0] io_right_bits_8,
  input  [15:0] io_right_bits_9,
  input  [15:0] io_right_bits_10,
  input  [15:0] io_right_bits_11,
  input  [15:0] io_right_bits_12,
  input  [15:0] io_right_bits_13,
  input  [15:0] io_right_bits_14,
  input  [15:0] io_right_bits_15,
  input  [15:0] io_right_bits_16,
  input  [15:0] io_right_bits_17,
  input  [15:0] io_right_bits_18,
  input  [15:0] io_right_bits_19,
  input  [15:0] io_right_bits_20,
  input  [15:0] io_right_bits_21,
  input  [15:0] io_right_bits_22,
  input  [15:0] io_right_bits_23,
  input  [15:0] io_right_bits_24,
  input  [15:0] io_right_bits_25,
  input  [15:0] io_right_bits_26,
  input  [15:0] io_right_bits_27,
  input  [15:0] io_right_bits_28,
  input  [15:0] io_right_bits_29,
  input  [15:0] io_right_bits_30,
  input  [15:0] io_right_bits_31,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_0,
  output [15:0] io_output_bits_1,
  output [15:0] io_output_bits_2,
  output [15:0] io_output_bits_3,
  output [15:0] io_output_bits_4,
  output [15:0] io_output_bits_5,
  output [15:0] io_output_bits_6,
  output [15:0] io_output_bits_7,
  output [15:0] io_output_bits_8,
  output [15:0] io_output_bits_9,
  output [15:0] io_output_bits_10,
  output [15:0] io_output_bits_11,
  output [15:0] io_output_bits_12,
  output [15:0] io_output_bits_13,
  output [15:0] io_output_bits_14,
  output [15:0] io_output_bits_15,
  output [15:0] io_output_bits_16,
  output [15:0] io_output_bits_17,
  output [15:0] io_output_bits_18,
  output [15:0] io_output_bits_19,
  output [15:0] io_output_bits_20,
  output [15:0] io_output_bits_21,
  output [15:0] io_output_bits_22,
  output [15:0] io_output_bits_23,
  output [15:0] io_output_bits_24,
  output [15:0] io_output_bits_25,
  output [15:0] io_output_bits_26,
  output [15:0] io_output_bits_27,
  output [15:0] io_output_bits_28,
  output [15:0] io_output_bits_29,
  output [15:0] io_output_bits_30,
  output [15:0] io_output_bits_31
);
  wire [25:0] _io_output_bits_0_mac_T = $signed(io_left_bits_0) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_0_mac_T_1 = {$signed(io_right_bits_0), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_0 = {{2{_io_output_bits_0_mac_T_1[23]}},_io_output_bits_0_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_0_mac = $signed(_io_output_bits_0_mac_T) + $signed(_GEN_0); // @[package.scala 117:23]
  wire [8:0] io_output_bits_0_mask1 = 9'sh80 - 9'sh1; // @[package.scala 120:44]
  wire [26:0] _io_output_bits_0_adjustment_T_1 = $signed(io_output_bits_0_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _GEN_1 = {{18{io_output_bits_0_mask1[8]}},io_output_bits_0_mask1}; // @[package.scala 125:44]
  wire [26:0] _io_output_bits_0_adjustment_T_4 = $signed(io_output_bits_0_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_0_adjustment_T_7 = $signed(io_output_bits_0_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_0_adjustment_T_10 = $signed(_io_output_bits_0_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_0_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_0_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_0_adjustment = _io_output_bits_0_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_0_adjusted_T = io_output_bits_0_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_2 = {{17{io_output_bits_0_adjustment[1]}},io_output_bits_0_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_0_adjusted = $signed(_io_output_bits_0_adjusted_T) + $signed(_GEN_2); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_0_saturated_T_2 = $signed(io_output_bits_0_adjusted) < -19'sh8000 ? $signed(-19'sh8000) :
    $signed(io_output_bits_0_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_0_saturated = $signed(io_output_bits_0_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_0_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_1_mac_T = $signed(io_left_bits_1) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_1_mac_T_1 = {$signed(io_right_bits_1), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_3 = {{2{_io_output_bits_1_mac_T_1[23]}},_io_output_bits_1_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_1_mac = $signed(_io_output_bits_1_mac_T) + $signed(_GEN_3); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_1_adjustment_T_1 = $signed(io_output_bits_1_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_1_adjustment_T_4 = $signed(io_output_bits_1_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_1_adjustment_T_7 = $signed(io_output_bits_1_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_1_adjustment_T_10 = $signed(_io_output_bits_1_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_1_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_1_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_1_adjustment = _io_output_bits_1_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_1_adjusted_T = io_output_bits_1_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_5 = {{17{io_output_bits_1_adjustment[1]}},io_output_bits_1_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_1_adjusted = $signed(_io_output_bits_1_adjusted_T) + $signed(_GEN_5); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_1_saturated_T_2 = $signed(io_output_bits_1_adjusted) < -19'sh8000 ? $signed(-19'sh8000) :
    $signed(io_output_bits_1_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_1_saturated = $signed(io_output_bits_1_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_1_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_2_mac_T = $signed(io_left_bits_2) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_2_mac_T_1 = {$signed(io_right_bits_2), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_6 = {{2{_io_output_bits_2_mac_T_1[23]}},_io_output_bits_2_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_2_mac = $signed(_io_output_bits_2_mac_T) + $signed(_GEN_6); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_2_adjustment_T_1 = $signed(io_output_bits_2_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_2_adjustment_T_4 = $signed(io_output_bits_2_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_2_adjustment_T_7 = $signed(io_output_bits_2_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_2_adjustment_T_10 = $signed(_io_output_bits_2_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_2_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_2_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_2_adjustment = _io_output_bits_2_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_2_adjusted_T = io_output_bits_2_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_8 = {{17{io_output_bits_2_adjustment[1]}},io_output_bits_2_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_2_adjusted = $signed(_io_output_bits_2_adjusted_T) + $signed(_GEN_8); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_2_saturated_T_2 = $signed(io_output_bits_2_adjusted) < -19'sh8000 ? $signed(-19'sh8000) :
    $signed(io_output_bits_2_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_2_saturated = $signed(io_output_bits_2_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_2_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_3_mac_T = $signed(io_left_bits_3) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_3_mac_T_1 = {$signed(io_right_bits_3), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_9 = {{2{_io_output_bits_3_mac_T_1[23]}},_io_output_bits_3_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_3_mac = $signed(_io_output_bits_3_mac_T) + $signed(_GEN_9); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_3_adjustment_T_1 = $signed(io_output_bits_3_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_3_adjustment_T_4 = $signed(io_output_bits_3_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_3_adjustment_T_7 = $signed(io_output_bits_3_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_3_adjustment_T_10 = $signed(_io_output_bits_3_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_3_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_3_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_3_adjustment = _io_output_bits_3_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_3_adjusted_T = io_output_bits_3_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_11 = {{17{io_output_bits_3_adjustment[1]}},io_output_bits_3_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_3_adjusted = $signed(_io_output_bits_3_adjusted_T) + $signed(_GEN_11); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_3_saturated_T_2 = $signed(io_output_bits_3_adjusted) < -19'sh8000 ? $signed(-19'sh8000) :
    $signed(io_output_bits_3_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_3_saturated = $signed(io_output_bits_3_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_3_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_4_mac_T = $signed(io_left_bits_4) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_4_mac_T_1 = {$signed(io_right_bits_4), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_12 = {{2{_io_output_bits_4_mac_T_1[23]}},_io_output_bits_4_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_4_mac = $signed(_io_output_bits_4_mac_T) + $signed(_GEN_12); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_4_adjustment_T_1 = $signed(io_output_bits_4_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_4_adjustment_T_4 = $signed(io_output_bits_4_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_4_adjustment_T_7 = $signed(io_output_bits_4_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_4_adjustment_T_10 = $signed(_io_output_bits_4_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_4_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_4_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_4_adjustment = _io_output_bits_4_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_4_adjusted_T = io_output_bits_4_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_14 = {{17{io_output_bits_4_adjustment[1]}},io_output_bits_4_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_4_adjusted = $signed(_io_output_bits_4_adjusted_T) + $signed(_GEN_14); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_4_saturated_T_2 = $signed(io_output_bits_4_adjusted) < -19'sh8000 ? $signed(-19'sh8000) :
    $signed(io_output_bits_4_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_4_saturated = $signed(io_output_bits_4_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_4_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_5_mac_T = $signed(io_left_bits_5) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_5_mac_T_1 = {$signed(io_right_bits_5), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_15 = {{2{_io_output_bits_5_mac_T_1[23]}},_io_output_bits_5_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_5_mac = $signed(_io_output_bits_5_mac_T) + $signed(_GEN_15); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_5_adjustment_T_1 = $signed(io_output_bits_5_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_5_adjustment_T_4 = $signed(io_output_bits_5_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_5_adjustment_T_7 = $signed(io_output_bits_5_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_5_adjustment_T_10 = $signed(_io_output_bits_5_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_5_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_5_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_5_adjustment = _io_output_bits_5_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_5_adjusted_T = io_output_bits_5_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_17 = {{17{io_output_bits_5_adjustment[1]}},io_output_bits_5_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_5_adjusted = $signed(_io_output_bits_5_adjusted_T) + $signed(_GEN_17); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_5_saturated_T_2 = $signed(io_output_bits_5_adjusted) < -19'sh8000 ? $signed(-19'sh8000) :
    $signed(io_output_bits_5_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_5_saturated = $signed(io_output_bits_5_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_5_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_6_mac_T = $signed(io_left_bits_6) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_6_mac_T_1 = {$signed(io_right_bits_6), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_18 = {{2{_io_output_bits_6_mac_T_1[23]}},_io_output_bits_6_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_6_mac = $signed(_io_output_bits_6_mac_T) + $signed(_GEN_18); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_6_adjustment_T_1 = $signed(io_output_bits_6_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_6_adjustment_T_4 = $signed(io_output_bits_6_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_6_adjustment_T_7 = $signed(io_output_bits_6_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_6_adjustment_T_10 = $signed(_io_output_bits_6_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_6_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_6_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_6_adjustment = _io_output_bits_6_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_6_adjusted_T = io_output_bits_6_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_20 = {{17{io_output_bits_6_adjustment[1]}},io_output_bits_6_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_6_adjusted = $signed(_io_output_bits_6_adjusted_T) + $signed(_GEN_20); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_6_saturated_T_2 = $signed(io_output_bits_6_adjusted) < -19'sh8000 ? $signed(-19'sh8000) :
    $signed(io_output_bits_6_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_6_saturated = $signed(io_output_bits_6_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_6_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_7_mac_T = $signed(io_left_bits_7) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_7_mac_T_1 = {$signed(io_right_bits_7), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_21 = {{2{_io_output_bits_7_mac_T_1[23]}},_io_output_bits_7_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_7_mac = $signed(_io_output_bits_7_mac_T) + $signed(_GEN_21); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_7_adjustment_T_1 = $signed(io_output_bits_7_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_7_adjustment_T_4 = $signed(io_output_bits_7_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_7_adjustment_T_7 = $signed(io_output_bits_7_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_7_adjustment_T_10 = $signed(_io_output_bits_7_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_7_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_7_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_7_adjustment = _io_output_bits_7_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_7_adjusted_T = io_output_bits_7_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_23 = {{17{io_output_bits_7_adjustment[1]}},io_output_bits_7_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_7_adjusted = $signed(_io_output_bits_7_adjusted_T) + $signed(_GEN_23); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_7_saturated_T_2 = $signed(io_output_bits_7_adjusted) < -19'sh8000 ? $signed(-19'sh8000) :
    $signed(io_output_bits_7_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_7_saturated = $signed(io_output_bits_7_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_7_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_8_mac_T = $signed(io_left_bits_8) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_8_mac_T_1 = {$signed(io_right_bits_8), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_24 = {{2{_io_output_bits_8_mac_T_1[23]}},_io_output_bits_8_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_8_mac = $signed(_io_output_bits_8_mac_T) + $signed(_GEN_24); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_8_adjustment_T_1 = $signed(io_output_bits_8_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_8_adjustment_T_4 = $signed(io_output_bits_8_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_8_adjustment_T_7 = $signed(io_output_bits_8_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_8_adjustment_T_10 = $signed(_io_output_bits_8_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_8_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_8_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_8_adjustment = _io_output_bits_8_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_8_adjusted_T = io_output_bits_8_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_26 = {{17{io_output_bits_8_adjustment[1]}},io_output_bits_8_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_8_adjusted = $signed(_io_output_bits_8_adjusted_T) + $signed(_GEN_26); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_8_saturated_T_2 = $signed(io_output_bits_8_adjusted) < -19'sh8000 ? $signed(-19'sh8000) :
    $signed(io_output_bits_8_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_8_saturated = $signed(io_output_bits_8_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_8_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_9_mac_T = $signed(io_left_bits_9) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_9_mac_T_1 = {$signed(io_right_bits_9), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_27 = {{2{_io_output_bits_9_mac_T_1[23]}},_io_output_bits_9_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_9_mac = $signed(_io_output_bits_9_mac_T) + $signed(_GEN_27); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_9_adjustment_T_1 = $signed(io_output_bits_9_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_9_adjustment_T_4 = $signed(io_output_bits_9_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_9_adjustment_T_7 = $signed(io_output_bits_9_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_9_adjustment_T_10 = $signed(_io_output_bits_9_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_9_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_9_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_9_adjustment = _io_output_bits_9_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_9_adjusted_T = io_output_bits_9_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_29 = {{17{io_output_bits_9_adjustment[1]}},io_output_bits_9_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_9_adjusted = $signed(_io_output_bits_9_adjusted_T) + $signed(_GEN_29); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_9_saturated_T_2 = $signed(io_output_bits_9_adjusted) < -19'sh8000 ? $signed(-19'sh8000) :
    $signed(io_output_bits_9_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_9_saturated = $signed(io_output_bits_9_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_9_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_10_mac_T = $signed(io_left_bits_10) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_10_mac_T_1 = {$signed(io_right_bits_10), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_30 = {{2{_io_output_bits_10_mac_T_1[23]}},_io_output_bits_10_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_10_mac = $signed(_io_output_bits_10_mac_T) + $signed(_GEN_30); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_10_adjustment_T_1 = $signed(io_output_bits_10_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_10_adjustment_T_4 = $signed(io_output_bits_10_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_10_adjustment_T_7 = $signed(io_output_bits_10_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_10_adjustment_T_10 = $signed(_io_output_bits_10_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_10_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_10_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_10_adjustment = _io_output_bits_10_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_10_adjusted_T = io_output_bits_10_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_32 = {{17{io_output_bits_10_adjustment[1]}},io_output_bits_10_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_10_adjusted = $signed(_io_output_bits_10_adjusted_T) + $signed(_GEN_32); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_10_saturated_T_2 = $signed(io_output_bits_10_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_10_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_10_saturated = $signed(io_output_bits_10_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_10_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_11_mac_T = $signed(io_left_bits_11) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_11_mac_T_1 = {$signed(io_right_bits_11), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_33 = {{2{_io_output_bits_11_mac_T_1[23]}},_io_output_bits_11_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_11_mac = $signed(_io_output_bits_11_mac_T) + $signed(_GEN_33); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_11_adjustment_T_1 = $signed(io_output_bits_11_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_11_adjustment_T_4 = $signed(io_output_bits_11_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_11_adjustment_T_7 = $signed(io_output_bits_11_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_11_adjustment_T_10 = $signed(_io_output_bits_11_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_11_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_11_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_11_adjustment = _io_output_bits_11_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_11_adjusted_T = io_output_bits_11_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_35 = {{17{io_output_bits_11_adjustment[1]}},io_output_bits_11_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_11_adjusted = $signed(_io_output_bits_11_adjusted_T) + $signed(_GEN_35); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_11_saturated_T_2 = $signed(io_output_bits_11_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_11_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_11_saturated = $signed(io_output_bits_11_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_11_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_12_mac_T = $signed(io_left_bits_12) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_12_mac_T_1 = {$signed(io_right_bits_12), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_36 = {{2{_io_output_bits_12_mac_T_1[23]}},_io_output_bits_12_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_12_mac = $signed(_io_output_bits_12_mac_T) + $signed(_GEN_36); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_12_adjustment_T_1 = $signed(io_output_bits_12_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_12_adjustment_T_4 = $signed(io_output_bits_12_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_12_adjustment_T_7 = $signed(io_output_bits_12_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_12_adjustment_T_10 = $signed(_io_output_bits_12_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_12_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_12_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_12_adjustment = _io_output_bits_12_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_12_adjusted_T = io_output_bits_12_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_38 = {{17{io_output_bits_12_adjustment[1]}},io_output_bits_12_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_12_adjusted = $signed(_io_output_bits_12_adjusted_T) + $signed(_GEN_38); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_12_saturated_T_2 = $signed(io_output_bits_12_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_12_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_12_saturated = $signed(io_output_bits_12_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_12_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_13_mac_T = $signed(io_left_bits_13) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_13_mac_T_1 = {$signed(io_right_bits_13), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_39 = {{2{_io_output_bits_13_mac_T_1[23]}},_io_output_bits_13_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_13_mac = $signed(_io_output_bits_13_mac_T) + $signed(_GEN_39); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_13_adjustment_T_1 = $signed(io_output_bits_13_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_13_adjustment_T_4 = $signed(io_output_bits_13_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_13_adjustment_T_7 = $signed(io_output_bits_13_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_13_adjustment_T_10 = $signed(_io_output_bits_13_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_13_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_13_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_13_adjustment = _io_output_bits_13_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_13_adjusted_T = io_output_bits_13_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_41 = {{17{io_output_bits_13_adjustment[1]}},io_output_bits_13_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_13_adjusted = $signed(_io_output_bits_13_adjusted_T) + $signed(_GEN_41); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_13_saturated_T_2 = $signed(io_output_bits_13_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_13_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_13_saturated = $signed(io_output_bits_13_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_13_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_14_mac_T = $signed(io_left_bits_14) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_14_mac_T_1 = {$signed(io_right_bits_14), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_42 = {{2{_io_output_bits_14_mac_T_1[23]}},_io_output_bits_14_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_14_mac = $signed(_io_output_bits_14_mac_T) + $signed(_GEN_42); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_14_adjustment_T_1 = $signed(io_output_bits_14_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_14_adjustment_T_4 = $signed(io_output_bits_14_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_14_adjustment_T_7 = $signed(io_output_bits_14_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_14_adjustment_T_10 = $signed(_io_output_bits_14_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_14_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_14_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_14_adjustment = _io_output_bits_14_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_14_adjusted_T = io_output_bits_14_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_44 = {{17{io_output_bits_14_adjustment[1]}},io_output_bits_14_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_14_adjusted = $signed(_io_output_bits_14_adjusted_T) + $signed(_GEN_44); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_14_saturated_T_2 = $signed(io_output_bits_14_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_14_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_14_saturated = $signed(io_output_bits_14_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_14_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_15_mac_T = $signed(io_left_bits_15) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_15_mac_T_1 = {$signed(io_right_bits_15), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_45 = {{2{_io_output_bits_15_mac_T_1[23]}},_io_output_bits_15_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_15_mac = $signed(_io_output_bits_15_mac_T) + $signed(_GEN_45); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_15_adjustment_T_1 = $signed(io_output_bits_15_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_15_adjustment_T_4 = $signed(io_output_bits_15_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_15_adjustment_T_7 = $signed(io_output_bits_15_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_15_adjustment_T_10 = $signed(_io_output_bits_15_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_15_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_15_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_15_adjustment = _io_output_bits_15_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_15_adjusted_T = io_output_bits_15_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_47 = {{17{io_output_bits_15_adjustment[1]}},io_output_bits_15_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_15_adjusted = $signed(_io_output_bits_15_adjusted_T) + $signed(_GEN_47); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_15_saturated_T_2 = $signed(io_output_bits_15_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_15_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_15_saturated = $signed(io_output_bits_15_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_15_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_16_mac_T = $signed(io_left_bits_16) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_16_mac_T_1 = {$signed(io_right_bits_16), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_48 = {{2{_io_output_bits_16_mac_T_1[23]}},_io_output_bits_16_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_16_mac = $signed(_io_output_bits_16_mac_T) + $signed(_GEN_48); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_16_adjustment_T_1 = $signed(io_output_bits_16_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_16_adjustment_T_4 = $signed(io_output_bits_16_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_16_adjustment_T_7 = $signed(io_output_bits_16_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_16_adjustment_T_10 = $signed(_io_output_bits_16_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_16_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_16_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_16_adjustment = _io_output_bits_16_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_16_adjusted_T = io_output_bits_16_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_50 = {{17{io_output_bits_16_adjustment[1]}},io_output_bits_16_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_16_adjusted = $signed(_io_output_bits_16_adjusted_T) + $signed(_GEN_50); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_16_saturated_T_2 = $signed(io_output_bits_16_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_16_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_16_saturated = $signed(io_output_bits_16_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_16_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_17_mac_T = $signed(io_left_bits_17) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_17_mac_T_1 = {$signed(io_right_bits_17), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_51 = {{2{_io_output_bits_17_mac_T_1[23]}},_io_output_bits_17_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_17_mac = $signed(_io_output_bits_17_mac_T) + $signed(_GEN_51); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_17_adjustment_T_1 = $signed(io_output_bits_17_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_17_adjustment_T_4 = $signed(io_output_bits_17_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_17_adjustment_T_7 = $signed(io_output_bits_17_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_17_adjustment_T_10 = $signed(_io_output_bits_17_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_17_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_17_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_17_adjustment = _io_output_bits_17_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_17_adjusted_T = io_output_bits_17_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_53 = {{17{io_output_bits_17_adjustment[1]}},io_output_bits_17_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_17_adjusted = $signed(_io_output_bits_17_adjusted_T) + $signed(_GEN_53); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_17_saturated_T_2 = $signed(io_output_bits_17_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_17_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_17_saturated = $signed(io_output_bits_17_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_17_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_18_mac_T = $signed(io_left_bits_18) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_18_mac_T_1 = {$signed(io_right_bits_18), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_54 = {{2{_io_output_bits_18_mac_T_1[23]}},_io_output_bits_18_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_18_mac = $signed(_io_output_bits_18_mac_T) + $signed(_GEN_54); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_18_adjustment_T_1 = $signed(io_output_bits_18_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_18_adjustment_T_4 = $signed(io_output_bits_18_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_18_adjustment_T_7 = $signed(io_output_bits_18_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_18_adjustment_T_10 = $signed(_io_output_bits_18_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_18_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_18_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_18_adjustment = _io_output_bits_18_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_18_adjusted_T = io_output_bits_18_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_56 = {{17{io_output_bits_18_adjustment[1]}},io_output_bits_18_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_18_adjusted = $signed(_io_output_bits_18_adjusted_T) + $signed(_GEN_56); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_18_saturated_T_2 = $signed(io_output_bits_18_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_18_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_18_saturated = $signed(io_output_bits_18_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_18_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_19_mac_T = $signed(io_left_bits_19) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_19_mac_T_1 = {$signed(io_right_bits_19), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_57 = {{2{_io_output_bits_19_mac_T_1[23]}},_io_output_bits_19_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_19_mac = $signed(_io_output_bits_19_mac_T) + $signed(_GEN_57); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_19_adjustment_T_1 = $signed(io_output_bits_19_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_19_adjustment_T_4 = $signed(io_output_bits_19_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_19_adjustment_T_7 = $signed(io_output_bits_19_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_19_adjustment_T_10 = $signed(_io_output_bits_19_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_19_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_19_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_19_adjustment = _io_output_bits_19_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_19_adjusted_T = io_output_bits_19_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_59 = {{17{io_output_bits_19_adjustment[1]}},io_output_bits_19_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_19_adjusted = $signed(_io_output_bits_19_adjusted_T) + $signed(_GEN_59); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_19_saturated_T_2 = $signed(io_output_bits_19_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_19_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_19_saturated = $signed(io_output_bits_19_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_19_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_20_mac_T = $signed(io_left_bits_20) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_20_mac_T_1 = {$signed(io_right_bits_20), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_60 = {{2{_io_output_bits_20_mac_T_1[23]}},_io_output_bits_20_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_20_mac = $signed(_io_output_bits_20_mac_T) + $signed(_GEN_60); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_20_adjustment_T_1 = $signed(io_output_bits_20_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_20_adjustment_T_4 = $signed(io_output_bits_20_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_20_adjustment_T_7 = $signed(io_output_bits_20_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_20_adjustment_T_10 = $signed(_io_output_bits_20_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_20_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_20_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_20_adjustment = _io_output_bits_20_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_20_adjusted_T = io_output_bits_20_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_62 = {{17{io_output_bits_20_adjustment[1]}},io_output_bits_20_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_20_adjusted = $signed(_io_output_bits_20_adjusted_T) + $signed(_GEN_62); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_20_saturated_T_2 = $signed(io_output_bits_20_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_20_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_20_saturated = $signed(io_output_bits_20_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_20_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_21_mac_T = $signed(io_left_bits_21) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_21_mac_T_1 = {$signed(io_right_bits_21), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_63 = {{2{_io_output_bits_21_mac_T_1[23]}},_io_output_bits_21_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_21_mac = $signed(_io_output_bits_21_mac_T) + $signed(_GEN_63); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_21_adjustment_T_1 = $signed(io_output_bits_21_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_21_adjustment_T_4 = $signed(io_output_bits_21_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_21_adjustment_T_7 = $signed(io_output_bits_21_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_21_adjustment_T_10 = $signed(_io_output_bits_21_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_21_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_21_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_21_adjustment = _io_output_bits_21_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_21_adjusted_T = io_output_bits_21_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_65 = {{17{io_output_bits_21_adjustment[1]}},io_output_bits_21_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_21_adjusted = $signed(_io_output_bits_21_adjusted_T) + $signed(_GEN_65); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_21_saturated_T_2 = $signed(io_output_bits_21_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_21_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_21_saturated = $signed(io_output_bits_21_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_21_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_22_mac_T = $signed(io_left_bits_22) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_22_mac_T_1 = {$signed(io_right_bits_22), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_66 = {{2{_io_output_bits_22_mac_T_1[23]}},_io_output_bits_22_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_22_mac = $signed(_io_output_bits_22_mac_T) + $signed(_GEN_66); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_22_adjustment_T_1 = $signed(io_output_bits_22_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_22_adjustment_T_4 = $signed(io_output_bits_22_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_22_adjustment_T_7 = $signed(io_output_bits_22_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_22_adjustment_T_10 = $signed(_io_output_bits_22_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_22_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_22_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_22_adjustment = _io_output_bits_22_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_22_adjusted_T = io_output_bits_22_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_68 = {{17{io_output_bits_22_adjustment[1]}},io_output_bits_22_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_22_adjusted = $signed(_io_output_bits_22_adjusted_T) + $signed(_GEN_68); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_22_saturated_T_2 = $signed(io_output_bits_22_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_22_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_22_saturated = $signed(io_output_bits_22_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_22_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_23_mac_T = $signed(io_left_bits_23) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_23_mac_T_1 = {$signed(io_right_bits_23), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_69 = {{2{_io_output_bits_23_mac_T_1[23]}},_io_output_bits_23_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_23_mac = $signed(_io_output_bits_23_mac_T) + $signed(_GEN_69); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_23_adjustment_T_1 = $signed(io_output_bits_23_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_23_adjustment_T_4 = $signed(io_output_bits_23_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_23_adjustment_T_7 = $signed(io_output_bits_23_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_23_adjustment_T_10 = $signed(_io_output_bits_23_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_23_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_23_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_23_adjustment = _io_output_bits_23_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_23_adjusted_T = io_output_bits_23_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_71 = {{17{io_output_bits_23_adjustment[1]}},io_output_bits_23_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_23_adjusted = $signed(_io_output_bits_23_adjusted_T) + $signed(_GEN_71); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_23_saturated_T_2 = $signed(io_output_bits_23_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_23_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_23_saturated = $signed(io_output_bits_23_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_23_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_24_mac_T = $signed(io_left_bits_24) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_24_mac_T_1 = {$signed(io_right_bits_24), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_72 = {{2{_io_output_bits_24_mac_T_1[23]}},_io_output_bits_24_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_24_mac = $signed(_io_output_bits_24_mac_T) + $signed(_GEN_72); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_24_adjustment_T_1 = $signed(io_output_bits_24_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_24_adjustment_T_4 = $signed(io_output_bits_24_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_24_adjustment_T_7 = $signed(io_output_bits_24_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_24_adjustment_T_10 = $signed(_io_output_bits_24_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_24_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_24_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_24_adjustment = _io_output_bits_24_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_24_adjusted_T = io_output_bits_24_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_74 = {{17{io_output_bits_24_adjustment[1]}},io_output_bits_24_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_24_adjusted = $signed(_io_output_bits_24_adjusted_T) + $signed(_GEN_74); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_24_saturated_T_2 = $signed(io_output_bits_24_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_24_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_24_saturated = $signed(io_output_bits_24_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_24_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_25_mac_T = $signed(io_left_bits_25) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_25_mac_T_1 = {$signed(io_right_bits_25), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_75 = {{2{_io_output_bits_25_mac_T_1[23]}},_io_output_bits_25_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_25_mac = $signed(_io_output_bits_25_mac_T) + $signed(_GEN_75); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_25_adjustment_T_1 = $signed(io_output_bits_25_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_25_adjustment_T_4 = $signed(io_output_bits_25_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_25_adjustment_T_7 = $signed(io_output_bits_25_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_25_adjustment_T_10 = $signed(_io_output_bits_25_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_25_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_25_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_25_adjustment = _io_output_bits_25_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_25_adjusted_T = io_output_bits_25_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_77 = {{17{io_output_bits_25_adjustment[1]}},io_output_bits_25_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_25_adjusted = $signed(_io_output_bits_25_adjusted_T) + $signed(_GEN_77); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_25_saturated_T_2 = $signed(io_output_bits_25_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_25_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_25_saturated = $signed(io_output_bits_25_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_25_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_26_mac_T = $signed(io_left_bits_26) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_26_mac_T_1 = {$signed(io_right_bits_26), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_78 = {{2{_io_output_bits_26_mac_T_1[23]}},_io_output_bits_26_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_26_mac = $signed(_io_output_bits_26_mac_T) + $signed(_GEN_78); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_26_adjustment_T_1 = $signed(io_output_bits_26_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_26_adjustment_T_4 = $signed(io_output_bits_26_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_26_adjustment_T_7 = $signed(io_output_bits_26_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_26_adjustment_T_10 = $signed(_io_output_bits_26_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_26_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_26_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_26_adjustment = _io_output_bits_26_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_26_adjusted_T = io_output_bits_26_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_80 = {{17{io_output_bits_26_adjustment[1]}},io_output_bits_26_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_26_adjusted = $signed(_io_output_bits_26_adjusted_T) + $signed(_GEN_80); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_26_saturated_T_2 = $signed(io_output_bits_26_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_26_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_26_saturated = $signed(io_output_bits_26_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_26_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_27_mac_T = $signed(io_left_bits_27) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_27_mac_T_1 = {$signed(io_right_bits_27), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_81 = {{2{_io_output_bits_27_mac_T_1[23]}},_io_output_bits_27_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_27_mac = $signed(_io_output_bits_27_mac_T) + $signed(_GEN_81); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_27_adjustment_T_1 = $signed(io_output_bits_27_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_27_adjustment_T_4 = $signed(io_output_bits_27_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_27_adjustment_T_7 = $signed(io_output_bits_27_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_27_adjustment_T_10 = $signed(_io_output_bits_27_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_27_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_27_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_27_adjustment = _io_output_bits_27_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_27_adjusted_T = io_output_bits_27_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_83 = {{17{io_output_bits_27_adjustment[1]}},io_output_bits_27_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_27_adjusted = $signed(_io_output_bits_27_adjusted_T) + $signed(_GEN_83); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_27_saturated_T_2 = $signed(io_output_bits_27_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_27_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_27_saturated = $signed(io_output_bits_27_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_27_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_28_mac_T = $signed(io_left_bits_28) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_28_mac_T_1 = {$signed(io_right_bits_28), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_84 = {{2{_io_output_bits_28_mac_T_1[23]}},_io_output_bits_28_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_28_mac = $signed(_io_output_bits_28_mac_T) + $signed(_GEN_84); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_28_adjustment_T_1 = $signed(io_output_bits_28_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_28_adjustment_T_4 = $signed(io_output_bits_28_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_28_adjustment_T_7 = $signed(io_output_bits_28_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_28_adjustment_T_10 = $signed(_io_output_bits_28_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_28_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_28_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_28_adjustment = _io_output_bits_28_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_28_adjusted_T = io_output_bits_28_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_86 = {{17{io_output_bits_28_adjustment[1]}},io_output_bits_28_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_28_adjusted = $signed(_io_output_bits_28_adjusted_T) + $signed(_GEN_86); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_28_saturated_T_2 = $signed(io_output_bits_28_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_28_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_28_saturated = $signed(io_output_bits_28_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_28_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_29_mac_T = $signed(io_left_bits_29) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_29_mac_T_1 = {$signed(io_right_bits_29), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_87 = {{2{_io_output_bits_29_mac_T_1[23]}},_io_output_bits_29_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_29_mac = $signed(_io_output_bits_29_mac_T) + $signed(_GEN_87); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_29_adjustment_T_1 = $signed(io_output_bits_29_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_29_adjustment_T_4 = $signed(io_output_bits_29_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_29_adjustment_T_7 = $signed(io_output_bits_29_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_29_adjustment_T_10 = $signed(_io_output_bits_29_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_29_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_29_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_29_adjustment = _io_output_bits_29_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_29_adjusted_T = io_output_bits_29_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_89 = {{17{io_output_bits_29_adjustment[1]}},io_output_bits_29_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_29_adjusted = $signed(_io_output_bits_29_adjusted_T) + $signed(_GEN_89); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_29_saturated_T_2 = $signed(io_output_bits_29_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_29_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_29_saturated = $signed(io_output_bits_29_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_29_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_30_mac_T = $signed(io_left_bits_30) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_30_mac_T_1 = {$signed(io_right_bits_30), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_90 = {{2{_io_output_bits_30_mac_T_1[23]}},_io_output_bits_30_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_30_mac = $signed(_io_output_bits_30_mac_T) + $signed(_GEN_90); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_30_adjustment_T_1 = $signed(io_output_bits_30_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_30_adjustment_T_4 = $signed(io_output_bits_30_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_30_adjustment_T_7 = $signed(io_output_bits_30_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_30_adjustment_T_10 = $signed(_io_output_bits_30_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_30_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_30_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_30_adjustment = _io_output_bits_30_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_30_adjusted_T = io_output_bits_30_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_92 = {{17{io_output_bits_30_adjustment[1]}},io_output_bits_30_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_30_adjusted = $signed(_io_output_bits_30_adjusted_T) + $signed(_GEN_92); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_30_saturated_T_2 = $signed(io_output_bits_30_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_30_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_30_saturated = $signed(io_output_bits_30_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_30_saturated_T_2); // @[package.scala 98:8]
  wire [25:0] _io_output_bits_31_mac_T = $signed(io_left_bits_31) * 10'sh100; // @[package.scala 117:18]
  wire [23:0] _io_output_bits_31_mac_T_1 = {$signed(io_right_bits_31), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_93 = {{2{_io_output_bits_31_mac_T_1[23]}},_io_output_bits_31_mac_T_1}; // @[package.scala 117:23]
  wire [26:0] io_output_bits_31_mac = $signed(_io_output_bits_31_mac_T) + $signed(_GEN_93); // @[package.scala 117:23]
  wire [26:0] _io_output_bits_31_adjustment_T_1 = $signed(io_output_bits_31_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _io_output_bits_31_adjustment_T_4 = $signed(io_output_bits_31_mac) & $signed(_GEN_1); // @[package.scala 125:44]
  wire [26:0] _io_output_bits_31_adjustment_T_7 = $signed(io_output_bits_31_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _io_output_bits_31_adjustment_T_10 = $signed(_io_output_bits_31_adjustment_T_1) != 27'sh0 & ($signed(
    _io_output_bits_31_adjustment_T_4) != 27'sh0 | $signed(_io_output_bits_31_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] io_output_bits_31_adjustment = _io_output_bits_31_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _io_output_bits_31_adjusted_T = io_output_bits_31_mac[26:8]; // @[package.scala 130:26]
  wire [18:0] _GEN_95 = {{17{io_output_bits_31_adjustment[1]}},io_output_bits_31_adjustment}; // @[package.scala 130:42]
  wire [18:0] io_output_bits_31_adjusted = $signed(_io_output_bits_31_adjusted_T) + $signed(_GEN_95); // @[package.scala 130:42]
  wire [18:0] _io_output_bits_31_saturated_T_2 = $signed(io_output_bits_31_adjusted) < -19'sh8000 ? $signed(-19'sh8000)
     : $signed(io_output_bits_31_adjusted); // @[package.scala 98:26]
  wire [18:0] io_output_bits_31_saturated = $signed(io_output_bits_31_adjusted) > 19'sh7fff ? $signed(19'sh7fff) :
    $signed(_io_output_bits_31_saturated_T_2); // @[package.scala 98:8]
  assign io_left_ready = io_output_ready & io_right_valid; // @[VecAdder.scala 24:33]
  assign io_right_ready = io_output_ready & io_left_valid; // @[VecAdder.scala 25:34]
  assign io_output_valid = io_left_valid & io_right_valid; // @[VecAdder.scala 23:33]
  assign io_output_bits_0 = io_output_bits_0_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_1 = io_output_bits_1_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_2 = io_output_bits_2_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_3 = io_output_bits_3_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_4 = io_output_bits_4_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_5 = io_output_bits_5_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_6 = io_output_bits_6_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_7 = io_output_bits_7_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_8 = io_output_bits_8_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_9 = io_output_bits_9_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_10 = io_output_bits_10_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_11 = io_output_bits_11_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_12 = io_output_bits_12_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_13 = io_output_bits_13_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_14 = io_output_bits_14_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_15 = io_output_bits_15_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_16 = io_output_bits_16_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_17 = io_output_bits_17_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_18 = io_output_bits_18_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_19 = io_output_bits_19_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_20 = io_output_bits_20_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_21 = io_output_bits_21_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_22 = io_output_bits_22_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_23 = io_output_bits_23_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_24 = io_output_bits_24_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_25 = io_output_bits_25_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_26 = io_output_bits_26_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_27 = io_output_bits_27_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_28 = io_output_bits_28_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_29 = io_output_bits_29_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_30 = io_output_bits_30_saturated[15:0]; // @[VecAdder.scala 21:23]
  assign io_output_bits_31 = io_output_bits_31_saturated[15:0]; // @[VecAdder.scala 21:23]
endmodule
module LockPool_1(
  input         clock,
  input         reset,
  output        io_actor_0_in_ready,
  input         io_actor_0_in_valid,
  input         io_actor_0_in_bits_write,
  input  [11:0] io_actor_0_in_bits_address,
  input  [11:0] io_actor_0_in_bits_size,
  input         io_actor_0_out_ready,
  output        io_actor_0_out_valid,
  output        io_actor_0_out_bits_write,
  output [11:0] io_actor_0_out_bits_address,
  output        io_actor_1_in_ready,
  input         io_actor_1_in_valid,
  input  [11:0] io_actor_1_in_bits_address,
  input         io_actor_1_out_ready,
  output        io_actor_1_out_valid,
  output [11:0] io_actor_1_out_bits_address,
  output        io_lock_ready,
  input         io_lock_valid,
  input  [11:0] io_lock_bits_cond_address
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  lock_0_cond_write; // @[LockPool.scala 55:21]
  reg [11:0] lock_0_cond_address; // @[LockPool.scala 55:21]
  reg  lock_0_held; // @[LockPool.scala 55:21]
  wire  _block_blocked_T_2 = io_lock_ready & io_lock_valid; // @[Decoupled.scala 50:35]
  wire  block_blocked_1 = lock_0_held | _block_blocked_T_2; // @[LockPool.scala 70:55]
  wire  _incomingObserved_T = io_actor_0_out_ready & io_actor_0_in_valid; // @[Decoupled.scala 50:35]
  wire  _incomingObserved_T_6 = io_actor_0_in_bits_write & io_actor_0_in_bits_address == io_lock_bits_cond_address &
    io_actor_0_in_bits_size == 12'h0; // @[MemControl.scala 59:56]
  wire  incomingObserved = io_lock_valid & _incomingObserved_T & _incomingObserved_T_6; // @[LockPool.scala 98:58]
  wire  _observed_T_5 = io_actor_0_in_bits_write == lock_0_cond_write & io_actor_0_in_bits_address ==
    lock_0_cond_address & io_actor_0_in_bits_size == 12'h0; // @[MemControl.scala 59:56]
  wire  observed = _incomingObserved_T & _observed_T_5; // @[LockPool.scala 107:37]
  wire  _GEN_32 = io_lock_valid | lock_0_cond_write; // @[LockPool.scala 86:29 89:14 55:21]
  wire [11:0] _GEN_33 = io_lock_valid ? io_lock_bits_cond_address : lock_0_cond_address; // @[LockPool.scala 86:29 89:14 55:21]
  wire  _GEN_45 = io_lock_valid | lock_0_held; // @[LockPool.scala 86:29 87:14 55:21]
  assign io_actor_0_in_ready = io_actor_0_out_ready; // @[LockPool.scala 139:40]
  assign io_actor_0_out_valid = io_actor_0_in_valid; // @[LockPool.scala 139:40]
  assign io_actor_0_out_bits_write = io_actor_0_in_bits_write; // @[LockPool.scala 139:40]
  assign io_actor_0_out_bits_address = io_actor_0_in_bits_address; // @[LockPool.scala 139:40]
  assign io_actor_1_in_ready = ~block_blocked_1 & io_actor_1_out_ready; // @[LockPool.scala 66:13 71:20 73:24]
  assign io_actor_1_out_valid = ~block_blocked_1 & io_actor_1_in_valid; // @[LockPool.scala 71:20 Decoupled.scala 72:20 LockPool.scala 73:24]
  assign io_actor_1_out_bits_address = io_actor_1_in_bits_address; // @[LockPool.scala 139:40]
  assign io_lock_ready = 1'h1; // @[LockPool.scala 104:24]
  always @(posedge clock) begin
    if (reset) begin // @[LockPool.scala 55:21]
      lock_0_cond_write <= 1'h0; // @[LockPool.scala 55:21]
    end else if (lock_0_held) begin // @[LockPool.scala 108:18]
      if (observed) begin // @[LockPool.scala 109:22]
        if (!(incomingObserved)) begin // @[LockPool.scala 111:34]
          lock_0_cond_write <= _GEN_32;
        end
      end else begin
        lock_0_cond_write <= _GEN_32;
      end
    end else if (~incomingObserved) begin // @[LockPool.scala 131:33]
      lock_0_cond_write <= _GEN_32;
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_0_cond_address <= 12'h0; // @[LockPool.scala 55:21]
    end else if (lock_0_held) begin // @[LockPool.scala 108:18]
      if (observed) begin // @[LockPool.scala 109:22]
        if (!(incomingObserved)) begin // @[LockPool.scala 111:34]
          lock_0_cond_address <= _GEN_33;
        end
      end else begin
        lock_0_cond_address <= _GEN_33;
      end
    end else if (~incomingObserved) begin // @[LockPool.scala 131:33]
      lock_0_cond_address <= _GEN_33;
    end
    if (reset) begin // @[LockPool.scala 55:21]
      lock_0_held <= 1'h0; // @[LockPool.scala 55:21]
    end else if (lock_0_held) begin // @[LockPool.scala 108:18]
      if (observed) begin // @[LockPool.scala 109:22]
        if (incomingObserved) begin // @[LockPool.scala 111:34]
          lock_0_held <= 1'h0; // @[LockPool.scala 93:12]
        end else begin
          lock_0_held <= io_lock_valid;
        end
      end else begin
        lock_0_held <= _GEN_45;
      end
    end else if (~incomingObserved) begin // @[LockPool.scala 131:33]
      lock_0_held <= _GEN_45;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lock_0_cond_write = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  lock_0_cond_address = _RAND_1[11:0];
  _RAND_2 = {1{`RANDOM}};
  lock_0_held = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_14(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_write,
  input  [11:0] io_enq_bits_address,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_write,
  output [11:0] io_deq_bits_address,
  output [11:0] io_deq_bits_size
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  ram_write [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_en; // @[Decoupled.scala 259:95]
  reg [11:0] ram_address [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [11:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [11:0] ram_address_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 259:95]
  reg [11:0] ram_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [11:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [11:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_11 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_11 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_write_io_deq_bits_MPORT_en = 1'h1;
  assign ram_write_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_write_io_deq_bits_MPORT_data = ram_write[ram_write_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_write_MPORT_data = io_enq_bits_write;
  assign ram_write_MPORT_addr = 1'h0;
  assign ram_write_MPORT_mask = 1'h1;
  assign ram_write_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = 1'h0;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = 12'h0;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_write = empty ? io_enq_bits_write : ram_write_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_address = empty ? io_enq_bits_address : ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? 12'h0 : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_write_MPORT_en & ram_write_MPORT_mask) begin
      ram_write[ram_write_MPORT_addr] <= ram_write_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_write[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_address[initvar] = _RAND_1[11:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[11:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Demux(
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_0,
  input  [15:0] io_in_bits_1,
  input  [15:0] io_in_bits_2,
  input  [15:0] io_in_bits_3,
  input  [15:0] io_in_bits_4,
  input  [15:0] io_in_bits_5,
  input  [15:0] io_in_bits_6,
  input  [15:0] io_in_bits_7,
  input  [15:0] io_in_bits_8,
  input  [15:0] io_in_bits_9,
  input  [15:0] io_in_bits_10,
  input  [15:0] io_in_bits_11,
  input  [15:0] io_in_bits_12,
  input  [15:0] io_in_bits_13,
  input  [15:0] io_in_bits_14,
  input  [15:0] io_in_bits_15,
  input  [15:0] io_in_bits_16,
  input  [15:0] io_in_bits_17,
  input  [15:0] io_in_bits_18,
  input  [15:0] io_in_bits_19,
  input  [15:0] io_in_bits_20,
  input  [15:0] io_in_bits_21,
  input  [15:0] io_in_bits_22,
  input  [15:0] io_in_bits_23,
  input  [15:0] io_in_bits_24,
  input  [15:0] io_in_bits_25,
  input  [15:0] io_in_bits_26,
  input  [15:0] io_in_bits_27,
  input  [15:0] io_in_bits_28,
  input  [15:0] io_in_bits_29,
  input  [15:0] io_in_bits_30,
  input  [15:0] io_in_bits_31,
  output        io_sel_ready,
  input         io_sel_valid,
  input         io_sel_bits,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [15:0] io_out_0_bits_0,
  output [15:0] io_out_0_bits_1,
  output [15:0] io_out_0_bits_2,
  output [15:0] io_out_0_bits_3,
  output [15:0] io_out_0_bits_4,
  output [15:0] io_out_0_bits_5,
  output [15:0] io_out_0_bits_6,
  output [15:0] io_out_0_bits_7,
  output [15:0] io_out_0_bits_8,
  output [15:0] io_out_0_bits_9,
  output [15:0] io_out_0_bits_10,
  output [15:0] io_out_0_bits_11,
  output [15:0] io_out_0_bits_12,
  output [15:0] io_out_0_bits_13,
  output [15:0] io_out_0_bits_14,
  output [15:0] io_out_0_bits_15,
  output [15:0] io_out_0_bits_16,
  output [15:0] io_out_0_bits_17,
  output [15:0] io_out_0_bits_18,
  output [15:0] io_out_0_bits_19,
  output [15:0] io_out_0_bits_20,
  output [15:0] io_out_0_bits_21,
  output [15:0] io_out_0_bits_22,
  output [15:0] io_out_0_bits_23,
  output [15:0] io_out_0_bits_24,
  output [15:0] io_out_0_bits_25,
  output [15:0] io_out_0_bits_26,
  output [15:0] io_out_0_bits_27,
  output [15:0] io_out_0_bits_28,
  output [15:0] io_out_0_bits_29,
  output [15:0] io_out_0_bits_30,
  output [15:0] io_out_0_bits_31,
  input         io_out_1_ready,
  output        io_out_1_valid,
  output [15:0] io_out_1_bits_0,
  output [15:0] io_out_1_bits_1,
  output [15:0] io_out_1_bits_2,
  output [15:0] io_out_1_bits_3,
  output [15:0] io_out_1_bits_4,
  output [15:0] io_out_1_bits_5,
  output [15:0] io_out_1_bits_6,
  output [15:0] io_out_1_bits_7,
  output [15:0] io_out_1_bits_8,
  output [15:0] io_out_1_bits_9,
  output [15:0] io_out_1_bits_10,
  output [15:0] io_out_1_bits_11,
  output [15:0] io_out_1_bits_12,
  output [15:0] io_out_1_bits_13,
  output [15:0] io_out_1_bits_14,
  output [15:0] io_out_1_bits_15,
  output [15:0] io_out_1_bits_16,
  output [15:0] io_out_1_bits_17,
  output [15:0] io_out_1_bits_18,
  output [15:0] io_out_1_bits_19,
  output [15:0] io_out_1_bits_20,
  output [15:0] io_out_1_bits_21,
  output [15:0] io_out_1_bits_22,
  output [15:0] io_out_1_bits_23,
  output [15:0] io_out_1_bits_24,
  output [15:0] io_out_1_bits_25,
  output [15:0] io_out_1_bits_26,
  output [15:0] io_out_1_bits_27,
  output [15:0] io_out_1_bits_28,
  output [15:0] io_out_1_bits_29,
  output [15:0] io_out_1_bits_30,
  output [15:0] io_out_1_bits_31
);
  wire  _GEN_67 = io_sel_bits ? io_out_1_ready : io_out_0_ready; // @[Demux.scala 34:{25,25}]
  assign io_in_ready = io_sel_valid & _GEN_67; // @[Demux.scala 35:25]
  assign io_sel_ready = io_in_valid & _GEN_67; // @[Demux.scala 34:25]
  assign io_out_0_valid = ~io_sel_bits & (io_sel_valid & io_in_valid); // @[Demux.scala 33:{13,13} 28:15]
  assign io_out_0_bits_0 = ~io_sel_bits ? $signed(io_in_bits_0) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_1 = ~io_sel_bits ? $signed(io_in_bits_1) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_2 = ~io_sel_bits ? $signed(io_in_bits_2) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_3 = ~io_sel_bits ? $signed(io_in_bits_3) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_4 = ~io_sel_bits ? $signed(io_in_bits_4) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_5 = ~io_sel_bits ? $signed(io_in_bits_5) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_6 = ~io_sel_bits ? $signed(io_in_bits_6) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_7 = ~io_sel_bits ? $signed(io_in_bits_7) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_8 = ~io_sel_bits ? $signed(io_in_bits_8) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_9 = ~io_sel_bits ? $signed(io_in_bits_9) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_10 = ~io_sel_bits ? $signed(io_in_bits_10) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_11 = ~io_sel_bits ? $signed(io_in_bits_11) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_12 = ~io_sel_bits ? $signed(io_in_bits_12) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_13 = ~io_sel_bits ? $signed(io_in_bits_13) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_14 = ~io_sel_bits ? $signed(io_in_bits_14) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_15 = ~io_sel_bits ? $signed(io_in_bits_15) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_16 = ~io_sel_bits ? $signed(io_in_bits_16) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_17 = ~io_sel_bits ? $signed(io_in_bits_17) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_18 = ~io_sel_bits ? $signed(io_in_bits_18) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_19 = ~io_sel_bits ? $signed(io_in_bits_19) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_20 = ~io_sel_bits ? $signed(io_in_bits_20) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_21 = ~io_sel_bits ? $signed(io_in_bits_21) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_22 = ~io_sel_bits ? $signed(io_in_bits_22) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_23 = ~io_sel_bits ? $signed(io_in_bits_23) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_24 = ~io_sel_bits ? $signed(io_in_bits_24) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_25 = ~io_sel_bits ? $signed(io_in_bits_25) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_26 = ~io_sel_bits ? $signed(io_in_bits_26) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_27 = ~io_sel_bits ? $signed(io_in_bits_27) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_28 = ~io_sel_bits ? $signed(io_in_bits_28) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_29 = ~io_sel_bits ? $signed(io_in_bits_29) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_30 = ~io_sel_bits ? $signed(io_in_bits_30) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_31 = ~io_sel_bits ? $signed(io_in_bits_31) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_valid = io_sel_bits & (io_sel_valid & io_in_valid); // @[Demux.scala 33:{13,13} 28:15]
  assign io_out_1_bits_0 = io_sel_bits ? $signed(io_in_bits_0) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_1 = io_sel_bits ? $signed(io_in_bits_1) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_2 = io_sel_bits ? $signed(io_in_bits_2) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_3 = io_sel_bits ? $signed(io_in_bits_3) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_4 = io_sel_bits ? $signed(io_in_bits_4) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_5 = io_sel_bits ? $signed(io_in_bits_5) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_6 = io_sel_bits ? $signed(io_in_bits_6) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_7 = io_sel_bits ? $signed(io_in_bits_7) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_8 = io_sel_bits ? $signed(io_in_bits_8) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_9 = io_sel_bits ? $signed(io_in_bits_9) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_10 = io_sel_bits ? $signed(io_in_bits_10) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_11 = io_sel_bits ? $signed(io_in_bits_11) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_12 = io_sel_bits ? $signed(io_in_bits_12) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_13 = io_sel_bits ? $signed(io_in_bits_13) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_14 = io_sel_bits ? $signed(io_in_bits_14) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_15 = io_sel_bits ? $signed(io_in_bits_15) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_16 = io_sel_bits ? $signed(io_in_bits_16) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_17 = io_sel_bits ? $signed(io_in_bits_17) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_18 = io_sel_bits ? $signed(io_in_bits_18) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_19 = io_sel_bits ? $signed(io_in_bits_19) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_20 = io_sel_bits ? $signed(io_in_bits_20) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_21 = io_sel_bits ? $signed(io_in_bits_21) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_22 = io_sel_bits ? $signed(io_in_bits_22) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_23 = io_sel_bits ? $signed(io_in_bits_23) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_24 = io_sel_bits ? $signed(io_in_bits_24) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_25 = io_sel_bits ? $signed(io_in_bits_25) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_26 = io_sel_bits ? $signed(io_in_bits_26) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_27 = io_sel_bits ? $signed(io_in_bits_27) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_28 = io_sel_bits ? $signed(io_in_bits_28) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_29 = io_sel_bits ? $signed(io_in_bits_29) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_30 = io_sel_bits ? $signed(io_in_bits_30) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_31 = io_sel_bits ? $signed(io_in_bits_31) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
endmodule
module Queue_15(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  ram [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_9 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_9 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = 1'h0;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = empty ? _GEN_9 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits = empty ? io_enq_bits : ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Mux(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [15:0] io_in_0_bits_0,
  input  [15:0] io_in_0_bits_1,
  input  [15:0] io_in_0_bits_2,
  input  [15:0] io_in_0_bits_3,
  input  [15:0] io_in_0_bits_4,
  input  [15:0] io_in_0_bits_5,
  input  [15:0] io_in_0_bits_6,
  input  [15:0] io_in_0_bits_7,
  input  [15:0] io_in_0_bits_8,
  input  [15:0] io_in_0_bits_9,
  input  [15:0] io_in_0_bits_10,
  input  [15:0] io_in_0_bits_11,
  input  [15:0] io_in_0_bits_12,
  input  [15:0] io_in_0_bits_13,
  input  [15:0] io_in_0_bits_14,
  input  [15:0] io_in_0_bits_15,
  input  [15:0] io_in_0_bits_16,
  input  [15:0] io_in_0_bits_17,
  input  [15:0] io_in_0_bits_18,
  input  [15:0] io_in_0_bits_19,
  input  [15:0] io_in_0_bits_20,
  input  [15:0] io_in_0_bits_21,
  input  [15:0] io_in_0_bits_22,
  input  [15:0] io_in_0_bits_23,
  input  [15:0] io_in_0_bits_24,
  input  [15:0] io_in_0_bits_25,
  input  [15:0] io_in_0_bits_26,
  input  [15:0] io_in_0_bits_27,
  input  [15:0] io_in_0_bits_28,
  input  [15:0] io_in_0_bits_29,
  input  [15:0] io_in_0_bits_30,
  input  [15:0] io_in_0_bits_31,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [15:0] io_in_1_bits_0,
  input  [15:0] io_in_1_bits_1,
  input  [15:0] io_in_1_bits_2,
  input  [15:0] io_in_1_bits_3,
  input  [15:0] io_in_1_bits_4,
  input  [15:0] io_in_1_bits_5,
  input  [15:0] io_in_1_bits_6,
  input  [15:0] io_in_1_bits_7,
  input  [15:0] io_in_1_bits_8,
  input  [15:0] io_in_1_bits_9,
  input  [15:0] io_in_1_bits_10,
  input  [15:0] io_in_1_bits_11,
  input  [15:0] io_in_1_bits_12,
  input  [15:0] io_in_1_bits_13,
  input  [15:0] io_in_1_bits_14,
  input  [15:0] io_in_1_bits_15,
  input  [15:0] io_in_1_bits_16,
  input  [15:0] io_in_1_bits_17,
  input  [15:0] io_in_1_bits_18,
  input  [15:0] io_in_1_bits_19,
  input  [15:0] io_in_1_bits_20,
  input  [15:0] io_in_1_bits_21,
  input  [15:0] io_in_1_bits_22,
  input  [15:0] io_in_1_bits_23,
  input  [15:0] io_in_1_bits_24,
  input  [15:0] io_in_1_bits_25,
  input  [15:0] io_in_1_bits_26,
  input  [15:0] io_in_1_bits_27,
  input  [15:0] io_in_1_bits_28,
  input  [15:0] io_in_1_bits_29,
  input  [15:0] io_in_1_bits_30,
  input  [15:0] io_in_1_bits_31,
  output        io_sel_ready,
  input         io_sel_valid,
  input         io_sel_bits,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_0,
  output [15:0] io_out_bits_1,
  output [15:0] io_out_bits_2,
  output [15:0] io_out_bits_3,
  output [15:0] io_out_bits_4,
  output [15:0] io_out_bits_5,
  output [15:0] io_out_bits_6,
  output [15:0] io_out_bits_7,
  output [15:0] io_out_bits_8,
  output [15:0] io_out_bits_9,
  output [15:0] io_out_bits_10,
  output [15:0] io_out_bits_11,
  output [15:0] io_out_bits_12,
  output [15:0] io_out_bits_13,
  output [15:0] io_out_bits_14,
  output [15:0] io_out_bits_15,
  output [15:0] io_out_bits_16,
  output [15:0] io_out_bits_17,
  output [15:0] io_out_bits_18,
  output [15:0] io_out_bits_19,
  output [15:0] io_out_bits_20,
  output [15:0] io_out_bits_21,
  output [15:0] io_out_bits_22,
  output [15:0] io_out_bits_23,
  output [15:0] io_out_bits_24,
  output [15:0] io_out_bits_25,
  output [15:0] io_out_bits_26,
  output [15:0] io_out_bits_27,
  output [15:0] io_out_bits_28,
  output [15:0] io_out_bits_29,
  output [15:0] io_out_bits_30,
  output [15:0] io_out_bits_31
);
  wire  _GEN_65 = io_sel_bits ? io_in_1_valid : io_in_0_valid; // @[Mux.scala 58:{29,29}]
  assign io_in_0_ready = ~io_sel_bits & (io_sel_valid & io_out_ready); // @[Mux.scala 60:{13,13} 52:19]
  assign io_in_1_ready = io_sel_bits & (io_sel_valid & io_out_ready); // @[Mux.scala 60:{13,13} 52:19]
  assign io_sel_ready = _GEN_65 & io_out_ready; // @[Mux.scala 59:26]
  assign io_out_valid = io_sel_valid & _GEN_65; // @[Mux.scala 58:29]
  assign io_out_bits_0 = io_sel_bits ? $signed(io_in_1_bits_0) : $signed(io_in_0_bits_0); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_1 = io_sel_bits ? $signed(io_in_1_bits_1) : $signed(io_in_0_bits_1); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_2 = io_sel_bits ? $signed(io_in_1_bits_2) : $signed(io_in_0_bits_2); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_3 = io_sel_bits ? $signed(io_in_1_bits_3) : $signed(io_in_0_bits_3); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_4 = io_sel_bits ? $signed(io_in_1_bits_4) : $signed(io_in_0_bits_4); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_5 = io_sel_bits ? $signed(io_in_1_bits_5) : $signed(io_in_0_bits_5); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_6 = io_sel_bits ? $signed(io_in_1_bits_6) : $signed(io_in_0_bits_6); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_7 = io_sel_bits ? $signed(io_in_1_bits_7) : $signed(io_in_0_bits_7); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_8 = io_sel_bits ? $signed(io_in_1_bits_8) : $signed(io_in_0_bits_8); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_9 = io_sel_bits ? $signed(io_in_1_bits_9) : $signed(io_in_0_bits_9); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_10 = io_sel_bits ? $signed(io_in_1_bits_10) : $signed(io_in_0_bits_10); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_11 = io_sel_bits ? $signed(io_in_1_bits_11) : $signed(io_in_0_bits_11); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_12 = io_sel_bits ? $signed(io_in_1_bits_12) : $signed(io_in_0_bits_12); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_13 = io_sel_bits ? $signed(io_in_1_bits_13) : $signed(io_in_0_bits_13); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_14 = io_sel_bits ? $signed(io_in_1_bits_14) : $signed(io_in_0_bits_14); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_15 = io_sel_bits ? $signed(io_in_1_bits_15) : $signed(io_in_0_bits_15); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_16 = io_sel_bits ? $signed(io_in_1_bits_16) : $signed(io_in_0_bits_16); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_17 = io_sel_bits ? $signed(io_in_1_bits_17) : $signed(io_in_0_bits_17); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_18 = io_sel_bits ? $signed(io_in_1_bits_18) : $signed(io_in_0_bits_18); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_19 = io_sel_bits ? $signed(io_in_1_bits_19) : $signed(io_in_0_bits_19); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_20 = io_sel_bits ? $signed(io_in_1_bits_20) : $signed(io_in_0_bits_20); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_21 = io_sel_bits ? $signed(io_in_1_bits_21) : $signed(io_in_0_bits_21); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_22 = io_sel_bits ? $signed(io_in_1_bits_22) : $signed(io_in_0_bits_22); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_23 = io_sel_bits ? $signed(io_in_1_bits_23) : $signed(io_in_0_bits_23); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_24 = io_sel_bits ? $signed(io_in_1_bits_24) : $signed(io_in_0_bits_24); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_25 = io_sel_bits ? $signed(io_in_1_bits_25) : $signed(io_in_0_bits_25); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_26 = io_sel_bits ? $signed(io_in_1_bits_26) : $signed(io_in_0_bits_26); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_27 = io_sel_bits ? $signed(io_in_1_bits_27) : $signed(io_in_0_bits_27); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_28 = io_sel_bits ? $signed(io_in_1_bits_28) : $signed(io_in_0_bits_28); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_29 = io_sel_bits ? $signed(io_in_1_bits_29) : $signed(io_in_0_bits_29); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_30 = io_sel_bits ? $signed(io_in_1_bits_30) : $signed(io_in_0_bits_30); // @[Mux.scala 57:{15,15}]
  assign io_out_bits_31 = io_sel_bits ? $signed(io_in_1_bits_31) : $signed(io_in_0_bits_31); // @[Mux.scala 57:{15,15}]
endmodule
module Accumulator(
  input         clock,
  input         reset,
  output        io_input_ready,
  input         io_input_valid,
  input  [15:0] io_input_bits_0,
  input  [15:0] io_input_bits_1,
  input  [15:0] io_input_bits_2,
  input  [15:0] io_input_bits_3,
  input  [15:0] io_input_bits_4,
  input  [15:0] io_input_bits_5,
  input  [15:0] io_input_bits_6,
  input  [15:0] io_input_bits_7,
  input  [15:0] io_input_bits_8,
  input  [15:0] io_input_bits_9,
  input  [15:0] io_input_bits_10,
  input  [15:0] io_input_bits_11,
  input  [15:0] io_input_bits_12,
  input  [15:0] io_input_bits_13,
  input  [15:0] io_input_bits_14,
  input  [15:0] io_input_bits_15,
  input  [15:0] io_input_bits_16,
  input  [15:0] io_input_bits_17,
  input  [15:0] io_input_bits_18,
  input  [15:0] io_input_bits_19,
  input  [15:0] io_input_bits_20,
  input  [15:0] io_input_bits_21,
  input  [15:0] io_input_bits_22,
  input  [15:0] io_input_bits_23,
  input  [15:0] io_input_bits_24,
  input  [15:0] io_input_bits_25,
  input  [15:0] io_input_bits_26,
  input  [15:0] io_input_bits_27,
  input  [15:0] io_input_bits_28,
  input  [15:0] io_input_bits_29,
  input  [15:0] io_input_bits_30,
  input  [15:0] io_input_bits_31,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_0,
  output [15:0] io_output_bits_1,
  output [15:0] io_output_bits_2,
  output [15:0] io_output_bits_3,
  output [15:0] io_output_bits_4,
  output [15:0] io_output_bits_5,
  output [15:0] io_output_bits_6,
  output [15:0] io_output_bits_7,
  output [15:0] io_output_bits_8,
  output [15:0] io_output_bits_9,
  output [15:0] io_output_bits_10,
  output [15:0] io_output_bits_11,
  output [15:0] io_output_bits_12,
  output [15:0] io_output_bits_13,
  output [15:0] io_output_bits_14,
  output [15:0] io_output_bits_15,
  output [15:0] io_output_bits_16,
  output [15:0] io_output_bits_17,
  output [15:0] io_output_bits_18,
  output [15:0] io_output_bits_19,
  output [15:0] io_output_bits_20,
  output [15:0] io_output_bits_21,
  output [15:0] io_output_bits_22,
  output [15:0] io_output_bits_23,
  output [15:0] io_output_bits_24,
  output [15:0] io_output_bits_25,
  output [15:0] io_output_bits_26,
  output [15:0] io_output_bits_27,
  output [15:0] io_output_bits_28,
  output [15:0] io_output_bits_29,
  output [15:0] io_output_bits_30,
  output [15:0] io_output_bits_31,
  output        io_control_ready,
  input         io_control_valid,
  input  [11:0] io_control_bits_address,
  input         io_control_bits_accumulate,
  input         io_control_bits_write,
  input         io_tracepoint,
  input  [31:0] io_programCounter
);
  wire  mem_clock; // @[Accumulator.scala 40:19]
  wire  mem_reset; // @[Accumulator.scala 40:19]
  wire  mem_io_portA_control_ready; // @[Accumulator.scala 40:19]
  wire  mem_io_portA_control_valid; // @[Accumulator.scala 40:19]
  wire  mem_io_portA_control_bits_write; // @[Accumulator.scala 40:19]
  wire [11:0] mem_io_portA_control_bits_address; // @[Accumulator.scala 40:19]
  wire  mem_io_portA_input_ready; // @[Accumulator.scala 40:19]
  wire  mem_io_portA_input_valid; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_0; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_1; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_2; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_3; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_4; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_5; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_6; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_7; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_8; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_9; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_10; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_11; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_12; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_13; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_14; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_15; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_16; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_17; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_18; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_19; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_20; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_21; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_22; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_23; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_24; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_25; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_26; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_27; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_28; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_29; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_30; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_input_bits_31; // @[Accumulator.scala 40:19]
  wire  mem_io_portA_output_ready; // @[Accumulator.scala 40:19]
  wire  mem_io_portA_output_valid; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_0; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_1; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_2; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_3; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_4; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_5; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_6; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_7; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_8; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_9; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_10; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_11; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_12; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_13; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_14; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_15; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_16; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_17; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_18; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_19; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_20; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_21; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_22; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_23; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_24; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_25; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_26; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_27; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_28; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_29; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_30; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portA_output_bits_31; // @[Accumulator.scala 40:19]
  wire  mem_io_portB_control_ready; // @[Accumulator.scala 40:19]
  wire  mem_io_portB_control_valid; // @[Accumulator.scala 40:19]
  wire [11:0] mem_io_portB_control_bits_address; // @[Accumulator.scala 40:19]
  wire  mem_io_portB_output_ready; // @[Accumulator.scala 40:19]
  wire  mem_io_portB_output_valid; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_0; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_1; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_2; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_3; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_4; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_5; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_6; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_7; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_8; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_9; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_10; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_11; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_12; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_13; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_14; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_15; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_16; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_17; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_18; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_19; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_20; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_21; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_22; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_23; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_24; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_25; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_26; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_27; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_28; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_29; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_30; // @[Accumulator.scala 40:19]
  wire [15:0] mem_io_portB_output_bits_31; // @[Accumulator.scala 40:19]
  wire  mem_io_tracepoint; // @[Accumulator.scala 40:19]
  wire [31:0] mem_io_programCounter; // @[Accumulator.scala 40:19]
  wire  adder_io_left_ready; // @[Accumulator.scala 49:23]
  wire  adder_io_left_valid; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_0; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_1; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_2; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_3; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_4; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_5; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_6; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_7; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_8; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_9; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_10; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_11; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_12; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_13; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_14; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_15; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_16; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_17; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_18; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_19; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_20; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_21; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_22; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_23; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_24; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_25; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_26; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_27; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_28; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_29; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_30; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_left_bits_31; // @[Accumulator.scala 49:23]
  wire  adder_io_right_ready; // @[Accumulator.scala 49:23]
  wire  adder_io_right_valid; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_0; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_1; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_2; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_3; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_4; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_5; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_6; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_7; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_8; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_9; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_10; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_11; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_12; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_13; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_14; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_15; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_16; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_17; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_18; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_19; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_20; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_21; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_22; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_23; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_24; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_25; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_26; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_27; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_28; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_29; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_30; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_right_bits_31; // @[Accumulator.scala 49:23]
  wire  adder_io_output_ready; // @[Accumulator.scala 49:23]
  wire  adder_io_output_valid; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_0; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_1; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_2; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_3; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_4; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_5; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_6; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_7; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_8; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_9; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_10; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_11; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_12; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_13; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_14; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_15; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_16; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_17; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_18; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_19; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_20; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_21; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_22; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_23; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_24; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_25; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_26; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_27; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_28; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_29; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_30; // @[Accumulator.scala 49:23]
  wire [15:0] adder_io_output_bits_31; // @[Accumulator.scala 49:23]
  wire  lockPool_clock; // @[Accumulator.scala 60:24]
  wire  lockPool_reset; // @[Accumulator.scala 60:24]
  wire  lockPool_io_actor_0_in_ready; // @[Accumulator.scala 60:24]
  wire  lockPool_io_actor_0_in_valid; // @[Accumulator.scala 60:24]
  wire  lockPool_io_actor_0_in_bits_write; // @[Accumulator.scala 60:24]
  wire [11:0] lockPool_io_actor_0_in_bits_address; // @[Accumulator.scala 60:24]
  wire [11:0] lockPool_io_actor_0_in_bits_size; // @[Accumulator.scala 60:24]
  wire  lockPool_io_actor_0_out_ready; // @[Accumulator.scala 60:24]
  wire  lockPool_io_actor_0_out_valid; // @[Accumulator.scala 60:24]
  wire  lockPool_io_actor_0_out_bits_write; // @[Accumulator.scala 60:24]
  wire [11:0] lockPool_io_actor_0_out_bits_address; // @[Accumulator.scala 60:24]
  wire  lockPool_io_actor_1_in_ready; // @[Accumulator.scala 60:24]
  wire  lockPool_io_actor_1_in_valid; // @[Accumulator.scala 60:24]
  wire [11:0] lockPool_io_actor_1_in_bits_address; // @[Accumulator.scala 60:24]
  wire  lockPool_io_actor_1_out_ready; // @[Accumulator.scala 60:24]
  wire  lockPool_io_actor_1_out_valid; // @[Accumulator.scala 60:24]
  wire [11:0] lockPool_io_actor_1_out_bits_address; // @[Accumulator.scala 60:24]
  wire  lockPool_io_lock_ready; // @[Accumulator.scala 60:24]
  wire  lockPool_io_lock_valid; // @[Accumulator.scala 60:24]
  wire [11:0] lockPool_io_lock_bits_cond_address; // @[Accumulator.scala 60:24]
  wire  portAControl_clock; // @[Mem.scala 22:19]
  wire  portAControl_reset; // @[Mem.scala 22:19]
  wire  portAControl_io_enq_ready; // @[Mem.scala 22:19]
  wire  portAControl_io_enq_valid; // @[Mem.scala 22:19]
  wire  portAControl_io_enq_bits_write; // @[Mem.scala 22:19]
  wire [11:0] portAControl_io_enq_bits_address; // @[Mem.scala 22:19]
  wire  portAControl_io_deq_ready; // @[Mem.scala 22:19]
  wire  portAControl_io_deq_valid; // @[Mem.scala 22:19]
  wire  portAControl_io_deq_bits_write; // @[Mem.scala 22:19]
  wire [11:0] portAControl_io_deq_bits_address; // @[Mem.scala 22:19]
  wire [11:0] portAControl_io_deq_bits_size; // @[Mem.scala 22:19]
  wire  inputDemuxModule_io_in_ready; // @[Accumulator.scala 88:32]
  wire  inputDemuxModule_io_in_valid; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_0; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_1; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_2; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_3; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_4; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_5; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_6; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_7; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_8; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_9; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_10; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_11; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_12; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_13; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_14; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_15; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_16; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_17; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_18; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_19; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_20; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_21; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_22; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_23; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_24; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_25; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_26; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_27; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_28; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_29; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_30; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_in_bits_31; // @[Accumulator.scala 88:32]
  wire  inputDemuxModule_io_sel_ready; // @[Accumulator.scala 88:32]
  wire  inputDemuxModule_io_sel_valid; // @[Accumulator.scala 88:32]
  wire  inputDemuxModule_io_sel_bits; // @[Accumulator.scala 88:32]
  wire  inputDemuxModule_io_out_0_ready; // @[Accumulator.scala 88:32]
  wire  inputDemuxModule_io_out_0_valid; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_0; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_1; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_2; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_3; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_4; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_5; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_6; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_7; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_8; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_9; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_10; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_11; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_12; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_13; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_14; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_15; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_16; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_17; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_18; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_19; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_20; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_21; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_22; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_23; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_24; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_25; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_26; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_27; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_28; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_29; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_30; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_0_bits_31; // @[Accumulator.scala 88:32]
  wire  inputDemuxModule_io_out_1_ready; // @[Accumulator.scala 88:32]
  wire  inputDemuxModule_io_out_1_valid; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_0; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_1; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_2; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_3; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_4; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_5; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_6; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_7; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_8; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_9; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_10; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_11; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_12; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_13; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_14; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_15; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_16; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_17; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_18; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_19; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_20; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_21; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_22; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_23; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_24; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_25; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_26; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_27; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_28; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_29; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_30; // @[Accumulator.scala 88:32]
  wire [15:0] inputDemuxModule_io_out_1_bits_31; // @[Accumulator.scala 88:32]
  wire  inputDemux_clock; // @[Mem.scala 22:19]
  wire  inputDemux_reset; // @[Mem.scala 22:19]
  wire  inputDemux_io_enq_ready; // @[Mem.scala 22:19]
  wire  inputDemux_io_enq_valid; // @[Mem.scala 22:19]
  wire  inputDemux_io_enq_bits; // @[Mem.scala 22:19]
  wire  inputDemux_io_deq_ready; // @[Mem.scala 22:19]
  wire  inputDemux_io_deq_valid; // @[Mem.scala 22:19]
  wire  inputDemux_io_deq_bits; // @[Mem.scala 22:19]
  wire  portAInputMux_x14_mux_io_in_0_ready; // @[Mux.scala 71:21]
  wire  portAInputMux_x14_mux_io_in_0_valid; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_0; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_1; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_2; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_3; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_4; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_5; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_6; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_7; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_8; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_9; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_10; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_11; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_12; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_13; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_14; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_15; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_16; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_17; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_18; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_19; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_20; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_21; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_22; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_23; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_24; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_25; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_26; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_27; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_28; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_29; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_30; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_0_bits_31; // @[Mux.scala 71:21]
  wire  portAInputMux_x14_mux_io_in_1_ready; // @[Mux.scala 71:21]
  wire  portAInputMux_x14_mux_io_in_1_valid; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_0; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_1; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_2; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_3; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_4; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_5; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_6; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_7; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_8; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_9; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_10; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_11; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_12; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_13; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_14; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_15; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_16; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_17; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_18; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_19; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_20; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_21; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_22; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_23; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_24; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_25; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_26; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_27; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_28; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_29; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_30; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_in_1_bits_31; // @[Mux.scala 71:21]
  wire  portAInputMux_x14_mux_io_sel_ready; // @[Mux.scala 71:21]
  wire  portAInputMux_x14_mux_io_sel_valid; // @[Mux.scala 71:21]
  wire  portAInputMux_x14_mux_io_sel_bits; // @[Mux.scala 71:21]
  wire  portAInputMux_x14_mux_io_out_ready; // @[Mux.scala 71:21]
  wire  portAInputMux_x14_mux_io_out_valid; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_0; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_1; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_2; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_3; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_4; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_5; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_6; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_7; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_8; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_9; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_10; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_11; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_12; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_13; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_14; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_15; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_16; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_17; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_18; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_19; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_20; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_21; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_22; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_23; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_24; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_25; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_26; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_27; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_28; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_29; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_30; // @[Mux.scala 71:21]
  wire [15:0] portAInputMux_x14_mux_io_out_bits_31; // @[Mux.scala 71:21]
  wire  portAInputMux_clock; // @[Mem.scala 22:19]
  wire  portAInputMux_reset; // @[Mem.scala 22:19]
  wire  portAInputMux_io_enq_ready; // @[Mem.scala 22:19]
  wire  portAInputMux_io_enq_valid; // @[Mem.scala 22:19]
  wire  portAInputMux_io_enq_bits; // @[Mem.scala 22:19]
  wire  portAInputMux_io_deq_ready; // @[Mem.scala 22:19]
  wire  portAInputMux_io_deq_valid; // @[Mem.scala 22:19]
  wire  portAInputMux_io_deq_bits; // @[Mem.scala 22:19]
  wire  writeEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_2_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_2_valid; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_3_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_3_valid; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_io_out_2_ready; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_io_out_2_valid; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_io_out_3_ready; // @[MultiEnqueue.scala 182:43]
  wire  accEnqueuer_io_out_3_valid; // @[MultiEnqueue.scala 182:43]
  wire  _GEN_0 = io_control_bits_accumulate & io_control_valid; // @[Accumulator.scala 112:35 MultiEnqueue.scala 150:17 40:17]
  wire  io_control_ready_portAControl_io_enq_w_ready = portAControl_io_enq_ready; // @[MultiEnqueue.scala 151:10 ReadyValid.scala 16:17]
  wire  _GEN_1 = io_control_bits_accumulate & io_control_ready_portAControl_io_enq_w_ready; // @[Accumulator.scala 112:35 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  io_control_ready_portAControl_io_enq_w_valid = accEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  io_control_ready_portAControl_io_enq_w_1_valid = writeEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_2 = io_control_bits_accumulate ? io_control_ready_portAControl_io_enq_w_valid :
    io_control_ready_portAControl_io_enq_w_1_valid; // @[Accumulator.scala 112:35 MultiEnqueue.scala 151:{10,10}]
  wire  io_control_ready_lockPool_io_actor_1_in_w_ready = lockPool_io_actor_1_in_ready; // @[MultiEnqueue.scala 152:10 ReadyValid.scala 16:17]
  wire  _GEN_6 = io_control_bits_accumulate & io_control_ready_lockPool_io_actor_1_in_w_ready; // @[Accumulator.scala 112:35 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  io_control_ready_lockPool_io_actor_1_in_w_valid = accEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_7 = io_control_bits_accumulate & io_control_ready_lockPool_io_actor_1_in_w_valid; // @[Accumulator.scala 112:35 MultiEnqueue.scala 152:10 package.scala 405:15]
  wire [11:0] _GEN_9 = io_control_bits_accumulate ? io_control_bits_address : 12'h0; // @[Accumulator.scala 112:35 MultiEnqueue.scala 152:10 package.scala 404:14]
  wire  io_control_ready_inputDemux_io_enq_w_ready = inputDemux_io_enq_ready; // @[MultiEnqueue.scala 153:10 ReadyValid.scala 16:17]
  wire  _GEN_11 = io_control_bits_accumulate & io_control_ready_inputDemux_io_enq_w_ready; // @[Accumulator.scala 112:35 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  io_control_ready_inputDemux_io_enq_w_valid = accEnqueuer_io_out_2_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  io_control_ready_inputDemux_io_enq_w_1_valid = writeEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_12 = io_control_bits_accumulate ? io_control_ready_inputDemux_io_enq_w_valid :
    io_control_ready_inputDemux_io_enq_w_1_valid; // @[Accumulator.scala 112:35 MultiEnqueue.scala 152:10 153:10]
  wire  io_control_ready_portAInputMux_io_enq_w_ready = portAInputMux_io_enq_ready; // @[MultiEnqueue.scala 154:10 ReadyValid.scala 16:17]
  wire  _GEN_14 = io_control_bits_accumulate & io_control_ready_portAInputMux_io_enq_w_ready; // @[Accumulator.scala 112:35 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  io_control_ready_portAInputMux_io_enq_w_valid = accEnqueuer_io_out_3_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  io_control_ready_portAInputMux_io_enq_w_1_valid = writeEnqueuer_io_out_2_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_15 = io_control_bits_accumulate ? io_control_ready_portAInputMux_io_enq_w_valid :
    io_control_ready_portAInputMux_io_enq_w_1_valid; // @[Accumulator.scala 112:35 MultiEnqueue.scala 153:10 154:10]
  wire  _GEN_17 = io_control_bits_accumulate ? accEnqueuer_io_in_ready : writeEnqueuer_io_in_ready; // @[Accumulator.scala 112:35 113:21 129:21]
  wire  _GEN_18 = io_control_bits_accumulate ? 1'h0 : io_control_valid; // @[Accumulator.scala 112:35 MultiEnqueue.scala 150:17 40:17]
  wire  _GEN_19 = io_control_bits_accumulate ? 1'h0 : io_control_ready_portAControl_io_enq_w_ready; // @[Accumulator.scala 112:35 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  _GEN_20 = io_control_bits_accumulate ? 1'h0 : io_control_ready_inputDemux_io_enq_w_ready; // @[Accumulator.scala 112:35 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  _GEN_21 = io_control_bits_accumulate ? 1'h0 : io_control_ready_portAInputMux_io_enq_w_ready; // @[Accumulator.scala 112:35 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  _GEN_22 = io_control_bits_accumulate ? 1'h0 : 1'h1; // @[Accumulator.scala 112:35 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  io_control_ready_lockPool_io_lock_w_valid = writeEnqueuer_io_out_3_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_23 = io_control_bits_accumulate ? 1'h0 : io_control_ready_lockPool_io_lock_w_valid; // @[Accumulator.scala 112:35 Decoupled.scala 72:20 MultiEnqueue.scala 154:10]
  wire  io_control_ready_portAControl_io_enq_w_2_valid = readEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  DualPortMem mem ( // @[Accumulator.scala 40:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_portA_control_ready(mem_io_portA_control_ready),
    .io_portA_control_valid(mem_io_portA_control_valid),
    .io_portA_control_bits_write(mem_io_portA_control_bits_write),
    .io_portA_control_bits_address(mem_io_portA_control_bits_address),
    .io_portA_input_ready(mem_io_portA_input_ready),
    .io_portA_input_valid(mem_io_portA_input_valid),
    .io_portA_input_bits_0(mem_io_portA_input_bits_0),
    .io_portA_input_bits_1(mem_io_portA_input_bits_1),
    .io_portA_input_bits_2(mem_io_portA_input_bits_2),
    .io_portA_input_bits_3(mem_io_portA_input_bits_3),
    .io_portA_input_bits_4(mem_io_portA_input_bits_4),
    .io_portA_input_bits_5(mem_io_portA_input_bits_5),
    .io_portA_input_bits_6(mem_io_portA_input_bits_6),
    .io_portA_input_bits_7(mem_io_portA_input_bits_7),
    .io_portA_input_bits_8(mem_io_portA_input_bits_8),
    .io_portA_input_bits_9(mem_io_portA_input_bits_9),
    .io_portA_input_bits_10(mem_io_portA_input_bits_10),
    .io_portA_input_bits_11(mem_io_portA_input_bits_11),
    .io_portA_input_bits_12(mem_io_portA_input_bits_12),
    .io_portA_input_bits_13(mem_io_portA_input_bits_13),
    .io_portA_input_bits_14(mem_io_portA_input_bits_14),
    .io_portA_input_bits_15(mem_io_portA_input_bits_15),
    .io_portA_input_bits_16(mem_io_portA_input_bits_16),
    .io_portA_input_bits_17(mem_io_portA_input_bits_17),
    .io_portA_input_bits_18(mem_io_portA_input_bits_18),
    .io_portA_input_bits_19(mem_io_portA_input_bits_19),
    .io_portA_input_bits_20(mem_io_portA_input_bits_20),
    .io_portA_input_bits_21(mem_io_portA_input_bits_21),
    .io_portA_input_bits_22(mem_io_portA_input_bits_22),
    .io_portA_input_bits_23(mem_io_portA_input_bits_23),
    .io_portA_input_bits_24(mem_io_portA_input_bits_24),
    .io_portA_input_bits_25(mem_io_portA_input_bits_25),
    .io_portA_input_bits_26(mem_io_portA_input_bits_26),
    .io_portA_input_bits_27(mem_io_portA_input_bits_27),
    .io_portA_input_bits_28(mem_io_portA_input_bits_28),
    .io_portA_input_bits_29(mem_io_portA_input_bits_29),
    .io_portA_input_bits_30(mem_io_portA_input_bits_30),
    .io_portA_input_bits_31(mem_io_portA_input_bits_31),
    .io_portA_output_ready(mem_io_portA_output_ready),
    .io_portA_output_valid(mem_io_portA_output_valid),
    .io_portA_output_bits_0(mem_io_portA_output_bits_0),
    .io_portA_output_bits_1(mem_io_portA_output_bits_1),
    .io_portA_output_bits_2(mem_io_portA_output_bits_2),
    .io_portA_output_bits_3(mem_io_portA_output_bits_3),
    .io_portA_output_bits_4(mem_io_portA_output_bits_4),
    .io_portA_output_bits_5(mem_io_portA_output_bits_5),
    .io_portA_output_bits_6(mem_io_portA_output_bits_6),
    .io_portA_output_bits_7(mem_io_portA_output_bits_7),
    .io_portA_output_bits_8(mem_io_portA_output_bits_8),
    .io_portA_output_bits_9(mem_io_portA_output_bits_9),
    .io_portA_output_bits_10(mem_io_portA_output_bits_10),
    .io_portA_output_bits_11(mem_io_portA_output_bits_11),
    .io_portA_output_bits_12(mem_io_portA_output_bits_12),
    .io_portA_output_bits_13(mem_io_portA_output_bits_13),
    .io_portA_output_bits_14(mem_io_portA_output_bits_14),
    .io_portA_output_bits_15(mem_io_portA_output_bits_15),
    .io_portA_output_bits_16(mem_io_portA_output_bits_16),
    .io_portA_output_bits_17(mem_io_portA_output_bits_17),
    .io_portA_output_bits_18(mem_io_portA_output_bits_18),
    .io_portA_output_bits_19(mem_io_portA_output_bits_19),
    .io_portA_output_bits_20(mem_io_portA_output_bits_20),
    .io_portA_output_bits_21(mem_io_portA_output_bits_21),
    .io_portA_output_bits_22(mem_io_portA_output_bits_22),
    .io_portA_output_bits_23(mem_io_portA_output_bits_23),
    .io_portA_output_bits_24(mem_io_portA_output_bits_24),
    .io_portA_output_bits_25(mem_io_portA_output_bits_25),
    .io_portA_output_bits_26(mem_io_portA_output_bits_26),
    .io_portA_output_bits_27(mem_io_portA_output_bits_27),
    .io_portA_output_bits_28(mem_io_portA_output_bits_28),
    .io_portA_output_bits_29(mem_io_portA_output_bits_29),
    .io_portA_output_bits_30(mem_io_portA_output_bits_30),
    .io_portA_output_bits_31(mem_io_portA_output_bits_31),
    .io_portB_control_ready(mem_io_portB_control_ready),
    .io_portB_control_valid(mem_io_portB_control_valid),
    .io_portB_control_bits_address(mem_io_portB_control_bits_address),
    .io_portB_output_ready(mem_io_portB_output_ready),
    .io_portB_output_valid(mem_io_portB_output_valid),
    .io_portB_output_bits_0(mem_io_portB_output_bits_0),
    .io_portB_output_bits_1(mem_io_portB_output_bits_1),
    .io_portB_output_bits_2(mem_io_portB_output_bits_2),
    .io_portB_output_bits_3(mem_io_portB_output_bits_3),
    .io_portB_output_bits_4(mem_io_portB_output_bits_4),
    .io_portB_output_bits_5(mem_io_portB_output_bits_5),
    .io_portB_output_bits_6(mem_io_portB_output_bits_6),
    .io_portB_output_bits_7(mem_io_portB_output_bits_7),
    .io_portB_output_bits_8(mem_io_portB_output_bits_8),
    .io_portB_output_bits_9(mem_io_portB_output_bits_9),
    .io_portB_output_bits_10(mem_io_portB_output_bits_10),
    .io_portB_output_bits_11(mem_io_portB_output_bits_11),
    .io_portB_output_bits_12(mem_io_portB_output_bits_12),
    .io_portB_output_bits_13(mem_io_portB_output_bits_13),
    .io_portB_output_bits_14(mem_io_portB_output_bits_14),
    .io_portB_output_bits_15(mem_io_portB_output_bits_15),
    .io_portB_output_bits_16(mem_io_portB_output_bits_16),
    .io_portB_output_bits_17(mem_io_portB_output_bits_17),
    .io_portB_output_bits_18(mem_io_portB_output_bits_18),
    .io_portB_output_bits_19(mem_io_portB_output_bits_19),
    .io_portB_output_bits_20(mem_io_portB_output_bits_20),
    .io_portB_output_bits_21(mem_io_portB_output_bits_21),
    .io_portB_output_bits_22(mem_io_portB_output_bits_22),
    .io_portB_output_bits_23(mem_io_portB_output_bits_23),
    .io_portB_output_bits_24(mem_io_portB_output_bits_24),
    .io_portB_output_bits_25(mem_io_portB_output_bits_25),
    .io_portB_output_bits_26(mem_io_portB_output_bits_26),
    .io_portB_output_bits_27(mem_io_portB_output_bits_27),
    .io_portB_output_bits_28(mem_io_portB_output_bits_28),
    .io_portB_output_bits_29(mem_io_portB_output_bits_29),
    .io_portB_output_bits_30(mem_io_portB_output_bits_30),
    .io_portB_output_bits_31(mem_io_portB_output_bits_31),
    .io_tracepoint(mem_io_tracepoint),
    .io_programCounter(mem_io_programCounter)
  );
  VecAdder adder ( // @[Accumulator.scala 49:23]
    .io_left_ready(adder_io_left_ready),
    .io_left_valid(adder_io_left_valid),
    .io_left_bits_0(adder_io_left_bits_0),
    .io_left_bits_1(adder_io_left_bits_1),
    .io_left_bits_2(adder_io_left_bits_2),
    .io_left_bits_3(adder_io_left_bits_3),
    .io_left_bits_4(adder_io_left_bits_4),
    .io_left_bits_5(adder_io_left_bits_5),
    .io_left_bits_6(adder_io_left_bits_6),
    .io_left_bits_7(adder_io_left_bits_7),
    .io_left_bits_8(adder_io_left_bits_8),
    .io_left_bits_9(adder_io_left_bits_9),
    .io_left_bits_10(adder_io_left_bits_10),
    .io_left_bits_11(adder_io_left_bits_11),
    .io_left_bits_12(adder_io_left_bits_12),
    .io_left_bits_13(adder_io_left_bits_13),
    .io_left_bits_14(adder_io_left_bits_14),
    .io_left_bits_15(adder_io_left_bits_15),
    .io_left_bits_16(adder_io_left_bits_16),
    .io_left_bits_17(adder_io_left_bits_17),
    .io_left_bits_18(adder_io_left_bits_18),
    .io_left_bits_19(adder_io_left_bits_19),
    .io_left_bits_20(adder_io_left_bits_20),
    .io_left_bits_21(adder_io_left_bits_21),
    .io_left_bits_22(adder_io_left_bits_22),
    .io_left_bits_23(adder_io_left_bits_23),
    .io_left_bits_24(adder_io_left_bits_24),
    .io_left_bits_25(adder_io_left_bits_25),
    .io_left_bits_26(adder_io_left_bits_26),
    .io_left_bits_27(adder_io_left_bits_27),
    .io_left_bits_28(adder_io_left_bits_28),
    .io_left_bits_29(adder_io_left_bits_29),
    .io_left_bits_30(adder_io_left_bits_30),
    .io_left_bits_31(adder_io_left_bits_31),
    .io_right_ready(adder_io_right_ready),
    .io_right_valid(adder_io_right_valid),
    .io_right_bits_0(adder_io_right_bits_0),
    .io_right_bits_1(adder_io_right_bits_1),
    .io_right_bits_2(adder_io_right_bits_2),
    .io_right_bits_3(adder_io_right_bits_3),
    .io_right_bits_4(adder_io_right_bits_4),
    .io_right_bits_5(adder_io_right_bits_5),
    .io_right_bits_6(adder_io_right_bits_6),
    .io_right_bits_7(adder_io_right_bits_7),
    .io_right_bits_8(adder_io_right_bits_8),
    .io_right_bits_9(adder_io_right_bits_9),
    .io_right_bits_10(adder_io_right_bits_10),
    .io_right_bits_11(adder_io_right_bits_11),
    .io_right_bits_12(adder_io_right_bits_12),
    .io_right_bits_13(adder_io_right_bits_13),
    .io_right_bits_14(adder_io_right_bits_14),
    .io_right_bits_15(adder_io_right_bits_15),
    .io_right_bits_16(adder_io_right_bits_16),
    .io_right_bits_17(adder_io_right_bits_17),
    .io_right_bits_18(adder_io_right_bits_18),
    .io_right_bits_19(adder_io_right_bits_19),
    .io_right_bits_20(adder_io_right_bits_20),
    .io_right_bits_21(adder_io_right_bits_21),
    .io_right_bits_22(adder_io_right_bits_22),
    .io_right_bits_23(adder_io_right_bits_23),
    .io_right_bits_24(adder_io_right_bits_24),
    .io_right_bits_25(adder_io_right_bits_25),
    .io_right_bits_26(adder_io_right_bits_26),
    .io_right_bits_27(adder_io_right_bits_27),
    .io_right_bits_28(adder_io_right_bits_28),
    .io_right_bits_29(adder_io_right_bits_29),
    .io_right_bits_30(adder_io_right_bits_30),
    .io_right_bits_31(adder_io_right_bits_31),
    .io_output_ready(adder_io_output_ready),
    .io_output_valid(adder_io_output_valid),
    .io_output_bits_0(adder_io_output_bits_0),
    .io_output_bits_1(adder_io_output_bits_1),
    .io_output_bits_2(adder_io_output_bits_2),
    .io_output_bits_3(adder_io_output_bits_3),
    .io_output_bits_4(adder_io_output_bits_4),
    .io_output_bits_5(adder_io_output_bits_5),
    .io_output_bits_6(adder_io_output_bits_6),
    .io_output_bits_7(adder_io_output_bits_7),
    .io_output_bits_8(adder_io_output_bits_8),
    .io_output_bits_9(adder_io_output_bits_9),
    .io_output_bits_10(adder_io_output_bits_10),
    .io_output_bits_11(adder_io_output_bits_11),
    .io_output_bits_12(adder_io_output_bits_12),
    .io_output_bits_13(adder_io_output_bits_13),
    .io_output_bits_14(adder_io_output_bits_14),
    .io_output_bits_15(adder_io_output_bits_15),
    .io_output_bits_16(adder_io_output_bits_16),
    .io_output_bits_17(adder_io_output_bits_17),
    .io_output_bits_18(adder_io_output_bits_18),
    .io_output_bits_19(adder_io_output_bits_19),
    .io_output_bits_20(adder_io_output_bits_20),
    .io_output_bits_21(adder_io_output_bits_21),
    .io_output_bits_22(adder_io_output_bits_22),
    .io_output_bits_23(adder_io_output_bits_23),
    .io_output_bits_24(adder_io_output_bits_24),
    .io_output_bits_25(adder_io_output_bits_25),
    .io_output_bits_26(adder_io_output_bits_26),
    .io_output_bits_27(adder_io_output_bits_27),
    .io_output_bits_28(adder_io_output_bits_28),
    .io_output_bits_29(adder_io_output_bits_29),
    .io_output_bits_30(adder_io_output_bits_30),
    .io_output_bits_31(adder_io_output_bits_31)
  );
  LockPool_1 lockPool ( // @[Accumulator.scala 60:24]
    .clock(lockPool_clock),
    .reset(lockPool_reset),
    .io_actor_0_in_ready(lockPool_io_actor_0_in_ready),
    .io_actor_0_in_valid(lockPool_io_actor_0_in_valid),
    .io_actor_0_in_bits_write(lockPool_io_actor_0_in_bits_write),
    .io_actor_0_in_bits_address(lockPool_io_actor_0_in_bits_address),
    .io_actor_0_in_bits_size(lockPool_io_actor_0_in_bits_size),
    .io_actor_0_out_ready(lockPool_io_actor_0_out_ready),
    .io_actor_0_out_valid(lockPool_io_actor_0_out_valid),
    .io_actor_0_out_bits_write(lockPool_io_actor_0_out_bits_write),
    .io_actor_0_out_bits_address(lockPool_io_actor_0_out_bits_address),
    .io_actor_1_in_ready(lockPool_io_actor_1_in_ready),
    .io_actor_1_in_valid(lockPool_io_actor_1_in_valid),
    .io_actor_1_in_bits_address(lockPool_io_actor_1_in_bits_address),
    .io_actor_1_out_ready(lockPool_io_actor_1_out_ready),
    .io_actor_1_out_valid(lockPool_io_actor_1_out_valid),
    .io_actor_1_out_bits_address(lockPool_io_actor_1_out_bits_address),
    .io_lock_ready(lockPool_io_lock_ready),
    .io_lock_valid(lockPool_io_lock_valid),
    .io_lock_bits_cond_address(lockPool_io_lock_bits_cond_address)
  );
  Queue_14 portAControl ( // @[Mem.scala 22:19]
    .clock(portAControl_clock),
    .reset(portAControl_reset),
    .io_enq_ready(portAControl_io_enq_ready),
    .io_enq_valid(portAControl_io_enq_valid),
    .io_enq_bits_write(portAControl_io_enq_bits_write),
    .io_enq_bits_address(portAControl_io_enq_bits_address),
    .io_deq_ready(portAControl_io_deq_ready),
    .io_deq_valid(portAControl_io_deq_valid),
    .io_deq_bits_write(portAControl_io_deq_bits_write),
    .io_deq_bits_address(portAControl_io_deq_bits_address),
    .io_deq_bits_size(portAControl_io_deq_bits_size)
  );
  Demux inputDemuxModule ( // @[Accumulator.scala 88:32]
    .io_in_ready(inputDemuxModule_io_in_ready),
    .io_in_valid(inputDemuxModule_io_in_valid),
    .io_in_bits_0(inputDemuxModule_io_in_bits_0),
    .io_in_bits_1(inputDemuxModule_io_in_bits_1),
    .io_in_bits_2(inputDemuxModule_io_in_bits_2),
    .io_in_bits_3(inputDemuxModule_io_in_bits_3),
    .io_in_bits_4(inputDemuxModule_io_in_bits_4),
    .io_in_bits_5(inputDemuxModule_io_in_bits_5),
    .io_in_bits_6(inputDemuxModule_io_in_bits_6),
    .io_in_bits_7(inputDemuxModule_io_in_bits_7),
    .io_in_bits_8(inputDemuxModule_io_in_bits_8),
    .io_in_bits_9(inputDemuxModule_io_in_bits_9),
    .io_in_bits_10(inputDemuxModule_io_in_bits_10),
    .io_in_bits_11(inputDemuxModule_io_in_bits_11),
    .io_in_bits_12(inputDemuxModule_io_in_bits_12),
    .io_in_bits_13(inputDemuxModule_io_in_bits_13),
    .io_in_bits_14(inputDemuxModule_io_in_bits_14),
    .io_in_bits_15(inputDemuxModule_io_in_bits_15),
    .io_in_bits_16(inputDemuxModule_io_in_bits_16),
    .io_in_bits_17(inputDemuxModule_io_in_bits_17),
    .io_in_bits_18(inputDemuxModule_io_in_bits_18),
    .io_in_bits_19(inputDemuxModule_io_in_bits_19),
    .io_in_bits_20(inputDemuxModule_io_in_bits_20),
    .io_in_bits_21(inputDemuxModule_io_in_bits_21),
    .io_in_bits_22(inputDemuxModule_io_in_bits_22),
    .io_in_bits_23(inputDemuxModule_io_in_bits_23),
    .io_in_bits_24(inputDemuxModule_io_in_bits_24),
    .io_in_bits_25(inputDemuxModule_io_in_bits_25),
    .io_in_bits_26(inputDemuxModule_io_in_bits_26),
    .io_in_bits_27(inputDemuxModule_io_in_bits_27),
    .io_in_bits_28(inputDemuxModule_io_in_bits_28),
    .io_in_bits_29(inputDemuxModule_io_in_bits_29),
    .io_in_bits_30(inputDemuxModule_io_in_bits_30),
    .io_in_bits_31(inputDemuxModule_io_in_bits_31),
    .io_sel_ready(inputDemuxModule_io_sel_ready),
    .io_sel_valid(inputDemuxModule_io_sel_valid),
    .io_sel_bits(inputDemuxModule_io_sel_bits),
    .io_out_0_ready(inputDemuxModule_io_out_0_ready),
    .io_out_0_valid(inputDemuxModule_io_out_0_valid),
    .io_out_0_bits_0(inputDemuxModule_io_out_0_bits_0),
    .io_out_0_bits_1(inputDemuxModule_io_out_0_bits_1),
    .io_out_0_bits_2(inputDemuxModule_io_out_0_bits_2),
    .io_out_0_bits_3(inputDemuxModule_io_out_0_bits_3),
    .io_out_0_bits_4(inputDemuxModule_io_out_0_bits_4),
    .io_out_0_bits_5(inputDemuxModule_io_out_0_bits_5),
    .io_out_0_bits_6(inputDemuxModule_io_out_0_bits_6),
    .io_out_0_bits_7(inputDemuxModule_io_out_0_bits_7),
    .io_out_0_bits_8(inputDemuxModule_io_out_0_bits_8),
    .io_out_0_bits_9(inputDemuxModule_io_out_0_bits_9),
    .io_out_0_bits_10(inputDemuxModule_io_out_0_bits_10),
    .io_out_0_bits_11(inputDemuxModule_io_out_0_bits_11),
    .io_out_0_bits_12(inputDemuxModule_io_out_0_bits_12),
    .io_out_0_bits_13(inputDemuxModule_io_out_0_bits_13),
    .io_out_0_bits_14(inputDemuxModule_io_out_0_bits_14),
    .io_out_0_bits_15(inputDemuxModule_io_out_0_bits_15),
    .io_out_0_bits_16(inputDemuxModule_io_out_0_bits_16),
    .io_out_0_bits_17(inputDemuxModule_io_out_0_bits_17),
    .io_out_0_bits_18(inputDemuxModule_io_out_0_bits_18),
    .io_out_0_bits_19(inputDemuxModule_io_out_0_bits_19),
    .io_out_0_bits_20(inputDemuxModule_io_out_0_bits_20),
    .io_out_0_bits_21(inputDemuxModule_io_out_0_bits_21),
    .io_out_0_bits_22(inputDemuxModule_io_out_0_bits_22),
    .io_out_0_bits_23(inputDemuxModule_io_out_0_bits_23),
    .io_out_0_bits_24(inputDemuxModule_io_out_0_bits_24),
    .io_out_0_bits_25(inputDemuxModule_io_out_0_bits_25),
    .io_out_0_bits_26(inputDemuxModule_io_out_0_bits_26),
    .io_out_0_bits_27(inputDemuxModule_io_out_0_bits_27),
    .io_out_0_bits_28(inputDemuxModule_io_out_0_bits_28),
    .io_out_0_bits_29(inputDemuxModule_io_out_0_bits_29),
    .io_out_0_bits_30(inputDemuxModule_io_out_0_bits_30),
    .io_out_0_bits_31(inputDemuxModule_io_out_0_bits_31),
    .io_out_1_ready(inputDemuxModule_io_out_1_ready),
    .io_out_1_valid(inputDemuxModule_io_out_1_valid),
    .io_out_1_bits_0(inputDemuxModule_io_out_1_bits_0),
    .io_out_1_bits_1(inputDemuxModule_io_out_1_bits_1),
    .io_out_1_bits_2(inputDemuxModule_io_out_1_bits_2),
    .io_out_1_bits_3(inputDemuxModule_io_out_1_bits_3),
    .io_out_1_bits_4(inputDemuxModule_io_out_1_bits_4),
    .io_out_1_bits_5(inputDemuxModule_io_out_1_bits_5),
    .io_out_1_bits_6(inputDemuxModule_io_out_1_bits_6),
    .io_out_1_bits_7(inputDemuxModule_io_out_1_bits_7),
    .io_out_1_bits_8(inputDemuxModule_io_out_1_bits_8),
    .io_out_1_bits_9(inputDemuxModule_io_out_1_bits_9),
    .io_out_1_bits_10(inputDemuxModule_io_out_1_bits_10),
    .io_out_1_bits_11(inputDemuxModule_io_out_1_bits_11),
    .io_out_1_bits_12(inputDemuxModule_io_out_1_bits_12),
    .io_out_1_bits_13(inputDemuxModule_io_out_1_bits_13),
    .io_out_1_bits_14(inputDemuxModule_io_out_1_bits_14),
    .io_out_1_bits_15(inputDemuxModule_io_out_1_bits_15),
    .io_out_1_bits_16(inputDemuxModule_io_out_1_bits_16),
    .io_out_1_bits_17(inputDemuxModule_io_out_1_bits_17),
    .io_out_1_bits_18(inputDemuxModule_io_out_1_bits_18),
    .io_out_1_bits_19(inputDemuxModule_io_out_1_bits_19),
    .io_out_1_bits_20(inputDemuxModule_io_out_1_bits_20),
    .io_out_1_bits_21(inputDemuxModule_io_out_1_bits_21),
    .io_out_1_bits_22(inputDemuxModule_io_out_1_bits_22),
    .io_out_1_bits_23(inputDemuxModule_io_out_1_bits_23),
    .io_out_1_bits_24(inputDemuxModule_io_out_1_bits_24),
    .io_out_1_bits_25(inputDemuxModule_io_out_1_bits_25),
    .io_out_1_bits_26(inputDemuxModule_io_out_1_bits_26),
    .io_out_1_bits_27(inputDemuxModule_io_out_1_bits_27),
    .io_out_1_bits_28(inputDemuxModule_io_out_1_bits_28),
    .io_out_1_bits_29(inputDemuxModule_io_out_1_bits_29),
    .io_out_1_bits_30(inputDemuxModule_io_out_1_bits_30),
    .io_out_1_bits_31(inputDemuxModule_io_out_1_bits_31)
  );
  Queue_15 inputDemux ( // @[Mem.scala 22:19]
    .clock(inputDemux_clock),
    .reset(inputDemux_reset),
    .io_enq_ready(inputDemux_io_enq_ready),
    .io_enq_valid(inputDemux_io_enq_valid),
    .io_enq_bits(inputDemux_io_enq_bits),
    .io_deq_ready(inputDemux_io_deq_ready),
    .io_deq_valid(inputDemux_io_deq_valid),
    .io_deq_bits(inputDemux_io_deq_bits)
  );
  Mux portAInputMux_x14_mux ( // @[Mux.scala 71:21]
    .io_in_0_ready(portAInputMux_x14_mux_io_in_0_ready),
    .io_in_0_valid(portAInputMux_x14_mux_io_in_0_valid),
    .io_in_0_bits_0(portAInputMux_x14_mux_io_in_0_bits_0),
    .io_in_0_bits_1(portAInputMux_x14_mux_io_in_0_bits_1),
    .io_in_0_bits_2(portAInputMux_x14_mux_io_in_0_bits_2),
    .io_in_0_bits_3(portAInputMux_x14_mux_io_in_0_bits_3),
    .io_in_0_bits_4(portAInputMux_x14_mux_io_in_0_bits_4),
    .io_in_0_bits_5(portAInputMux_x14_mux_io_in_0_bits_5),
    .io_in_0_bits_6(portAInputMux_x14_mux_io_in_0_bits_6),
    .io_in_0_bits_7(portAInputMux_x14_mux_io_in_0_bits_7),
    .io_in_0_bits_8(portAInputMux_x14_mux_io_in_0_bits_8),
    .io_in_0_bits_9(portAInputMux_x14_mux_io_in_0_bits_9),
    .io_in_0_bits_10(portAInputMux_x14_mux_io_in_0_bits_10),
    .io_in_0_bits_11(portAInputMux_x14_mux_io_in_0_bits_11),
    .io_in_0_bits_12(portAInputMux_x14_mux_io_in_0_bits_12),
    .io_in_0_bits_13(portAInputMux_x14_mux_io_in_0_bits_13),
    .io_in_0_bits_14(portAInputMux_x14_mux_io_in_0_bits_14),
    .io_in_0_bits_15(portAInputMux_x14_mux_io_in_0_bits_15),
    .io_in_0_bits_16(portAInputMux_x14_mux_io_in_0_bits_16),
    .io_in_0_bits_17(portAInputMux_x14_mux_io_in_0_bits_17),
    .io_in_0_bits_18(portAInputMux_x14_mux_io_in_0_bits_18),
    .io_in_0_bits_19(portAInputMux_x14_mux_io_in_0_bits_19),
    .io_in_0_bits_20(portAInputMux_x14_mux_io_in_0_bits_20),
    .io_in_0_bits_21(portAInputMux_x14_mux_io_in_0_bits_21),
    .io_in_0_bits_22(portAInputMux_x14_mux_io_in_0_bits_22),
    .io_in_0_bits_23(portAInputMux_x14_mux_io_in_0_bits_23),
    .io_in_0_bits_24(portAInputMux_x14_mux_io_in_0_bits_24),
    .io_in_0_bits_25(portAInputMux_x14_mux_io_in_0_bits_25),
    .io_in_0_bits_26(portAInputMux_x14_mux_io_in_0_bits_26),
    .io_in_0_bits_27(portAInputMux_x14_mux_io_in_0_bits_27),
    .io_in_0_bits_28(portAInputMux_x14_mux_io_in_0_bits_28),
    .io_in_0_bits_29(portAInputMux_x14_mux_io_in_0_bits_29),
    .io_in_0_bits_30(portAInputMux_x14_mux_io_in_0_bits_30),
    .io_in_0_bits_31(portAInputMux_x14_mux_io_in_0_bits_31),
    .io_in_1_ready(portAInputMux_x14_mux_io_in_1_ready),
    .io_in_1_valid(portAInputMux_x14_mux_io_in_1_valid),
    .io_in_1_bits_0(portAInputMux_x14_mux_io_in_1_bits_0),
    .io_in_1_bits_1(portAInputMux_x14_mux_io_in_1_bits_1),
    .io_in_1_bits_2(portAInputMux_x14_mux_io_in_1_bits_2),
    .io_in_1_bits_3(portAInputMux_x14_mux_io_in_1_bits_3),
    .io_in_1_bits_4(portAInputMux_x14_mux_io_in_1_bits_4),
    .io_in_1_bits_5(portAInputMux_x14_mux_io_in_1_bits_5),
    .io_in_1_bits_6(portAInputMux_x14_mux_io_in_1_bits_6),
    .io_in_1_bits_7(portAInputMux_x14_mux_io_in_1_bits_7),
    .io_in_1_bits_8(portAInputMux_x14_mux_io_in_1_bits_8),
    .io_in_1_bits_9(portAInputMux_x14_mux_io_in_1_bits_9),
    .io_in_1_bits_10(portAInputMux_x14_mux_io_in_1_bits_10),
    .io_in_1_bits_11(portAInputMux_x14_mux_io_in_1_bits_11),
    .io_in_1_bits_12(portAInputMux_x14_mux_io_in_1_bits_12),
    .io_in_1_bits_13(portAInputMux_x14_mux_io_in_1_bits_13),
    .io_in_1_bits_14(portAInputMux_x14_mux_io_in_1_bits_14),
    .io_in_1_bits_15(portAInputMux_x14_mux_io_in_1_bits_15),
    .io_in_1_bits_16(portAInputMux_x14_mux_io_in_1_bits_16),
    .io_in_1_bits_17(portAInputMux_x14_mux_io_in_1_bits_17),
    .io_in_1_bits_18(portAInputMux_x14_mux_io_in_1_bits_18),
    .io_in_1_bits_19(portAInputMux_x14_mux_io_in_1_bits_19),
    .io_in_1_bits_20(portAInputMux_x14_mux_io_in_1_bits_20),
    .io_in_1_bits_21(portAInputMux_x14_mux_io_in_1_bits_21),
    .io_in_1_bits_22(portAInputMux_x14_mux_io_in_1_bits_22),
    .io_in_1_bits_23(portAInputMux_x14_mux_io_in_1_bits_23),
    .io_in_1_bits_24(portAInputMux_x14_mux_io_in_1_bits_24),
    .io_in_1_bits_25(portAInputMux_x14_mux_io_in_1_bits_25),
    .io_in_1_bits_26(portAInputMux_x14_mux_io_in_1_bits_26),
    .io_in_1_bits_27(portAInputMux_x14_mux_io_in_1_bits_27),
    .io_in_1_bits_28(portAInputMux_x14_mux_io_in_1_bits_28),
    .io_in_1_bits_29(portAInputMux_x14_mux_io_in_1_bits_29),
    .io_in_1_bits_30(portAInputMux_x14_mux_io_in_1_bits_30),
    .io_in_1_bits_31(portAInputMux_x14_mux_io_in_1_bits_31),
    .io_sel_ready(portAInputMux_x14_mux_io_sel_ready),
    .io_sel_valid(portAInputMux_x14_mux_io_sel_valid),
    .io_sel_bits(portAInputMux_x14_mux_io_sel_bits),
    .io_out_ready(portAInputMux_x14_mux_io_out_ready),
    .io_out_valid(portAInputMux_x14_mux_io_out_valid),
    .io_out_bits_0(portAInputMux_x14_mux_io_out_bits_0),
    .io_out_bits_1(portAInputMux_x14_mux_io_out_bits_1),
    .io_out_bits_2(portAInputMux_x14_mux_io_out_bits_2),
    .io_out_bits_3(portAInputMux_x14_mux_io_out_bits_3),
    .io_out_bits_4(portAInputMux_x14_mux_io_out_bits_4),
    .io_out_bits_5(portAInputMux_x14_mux_io_out_bits_5),
    .io_out_bits_6(portAInputMux_x14_mux_io_out_bits_6),
    .io_out_bits_7(portAInputMux_x14_mux_io_out_bits_7),
    .io_out_bits_8(portAInputMux_x14_mux_io_out_bits_8),
    .io_out_bits_9(portAInputMux_x14_mux_io_out_bits_9),
    .io_out_bits_10(portAInputMux_x14_mux_io_out_bits_10),
    .io_out_bits_11(portAInputMux_x14_mux_io_out_bits_11),
    .io_out_bits_12(portAInputMux_x14_mux_io_out_bits_12),
    .io_out_bits_13(portAInputMux_x14_mux_io_out_bits_13),
    .io_out_bits_14(portAInputMux_x14_mux_io_out_bits_14),
    .io_out_bits_15(portAInputMux_x14_mux_io_out_bits_15),
    .io_out_bits_16(portAInputMux_x14_mux_io_out_bits_16),
    .io_out_bits_17(portAInputMux_x14_mux_io_out_bits_17),
    .io_out_bits_18(portAInputMux_x14_mux_io_out_bits_18),
    .io_out_bits_19(portAInputMux_x14_mux_io_out_bits_19),
    .io_out_bits_20(portAInputMux_x14_mux_io_out_bits_20),
    .io_out_bits_21(portAInputMux_x14_mux_io_out_bits_21),
    .io_out_bits_22(portAInputMux_x14_mux_io_out_bits_22),
    .io_out_bits_23(portAInputMux_x14_mux_io_out_bits_23),
    .io_out_bits_24(portAInputMux_x14_mux_io_out_bits_24),
    .io_out_bits_25(portAInputMux_x14_mux_io_out_bits_25),
    .io_out_bits_26(portAInputMux_x14_mux_io_out_bits_26),
    .io_out_bits_27(portAInputMux_x14_mux_io_out_bits_27),
    .io_out_bits_28(portAInputMux_x14_mux_io_out_bits_28),
    .io_out_bits_29(portAInputMux_x14_mux_io_out_bits_29),
    .io_out_bits_30(portAInputMux_x14_mux_io_out_bits_30),
    .io_out_bits_31(portAInputMux_x14_mux_io_out_bits_31)
  );
  Queue_15 portAInputMux ( // @[Mem.scala 22:19]
    .clock(portAInputMux_clock),
    .reset(portAInputMux_reset),
    .io_enq_ready(portAInputMux_io_enq_ready),
    .io_enq_valid(portAInputMux_io_enq_valid),
    .io_enq_bits(portAInputMux_io_enq_bits),
    .io_deq_ready(portAInputMux_io_deq_ready),
    .io_deq_valid(portAInputMux_io_deq_valid),
    .io_deq_bits(portAInputMux_io_deq_bits)
  );
  MultiEnqueue_3 writeEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(writeEnqueuer_clock),
    .reset(writeEnqueuer_reset),
    .io_in_ready(writeEnqueuer_io_in_ready),
    .io_in_valid(writeEnqueuer_io_in_valid),
    .io_out_0_ready(writeEnqueuer_io_out_0_ready),
    .io_out_0_valid(writeEnqueuer_io_out_0_valid),
    .io_out_1_ready(writeEnqueuer_io_out_1_ready),
    .io_out_1_valid(writeEnqueuer_io_out_1_valid),
    .io_out_2_ready(writeEnqueuer_io_out_2_ready),
    .io_out_2_valid(writeEnqueuer_io_out_2_valid),
    .io_out_3_ready(writeEnqueuer_io_out_3_ready),
    .io_out_3_valid(writeEnqueuer_io_out_3_valid)
  );
  MultiEnqueue readEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(readEnqueuer_clock),
    .reset(readEnqueuer_reset),
    .io_in_ready(readEnqueuer_io_in_ready),
    .io_in_valid(readEnqueuer_io_in_valid),
    .io_out_0_ready(readEnqueuer_io_out_0_ready),
    .io_out_0_valid(readEnqueuer_io_out_0_valid)
  );
  MultiEnqueue_3 accEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(accEnqueuer_clock),
    .reset(accEnqueuer_reset),
    .io_in_ready(accEnqueuer_io_in_ready),
    .io_in_valid(accEnqueuer_io_in_valid),
    .io_out_0_ready(accEnqueuer_io_out_0_ready),
    .io_out_0_valid(accEnqueuer_io_out_0_valid),
    .io_out_1_ready(accEnqueuer_io_out_1_ready),
    .io_out_1_valid(accEnqueuer_io_out_1_valid),
    .io_out_2_ready(accEnqueuer_io_out_2_ready),
    .io_out_2_valid(accEnqueuer_io_out_2_valid),
    .io_out_3_ready(accEnqueuer_io_out_3_ready),
    .io_out_3_valid(accEnqueuer_io_out_3_valid)
  );
  assign io_input_ready = inputDemuxModule_io_in_ready; // @[Accumulator.scala 93:26]
  assign io_output_valid = mem_io_portA_output_valid; // @[Accumulator.scala 84:13]
  assign io_output_bits_0 = mem_io_portA_output_bits_0; // @[Accumulator.scala 84:13]
  assign io_output_bits_1 = mem_io_portA_output_bits_1; // @[Accumulator.scala 84:13]
  assign io_output_bits_2 = mem_io_portA_output_bits_2; // @[Accumulator.scala 84:13]
  assign io_output_bits_3 = mem_io_portA_output_bits_3; // @[Accumulator.scala 84:13]
  assign io_output_bits_4 = mem_io_portA_output_bits_4; // @[Accumulator.scala 84:13]
  assign io_output_bits_5 = mem_io_portA_output_bits_5; // @[Accumulator.scala 84:13]
  assign io_output_bits_6 = mem_io_portA_output_bits_6; // @[Accumulator.scala 84:13]
  assign io_output_bits_7 = mem_io_portA_output_bits_7; // @[Accumulator.scala 84:13]
  assign io_output_bits_8 = mem_io_portA_output_bits_8; // @[Accumulator.scala 84:13]
  assign io_output_bits_9 = mem_io_portA_output_bits_9; // @[Accumulator.scala 84:13]
  assign io_output_bits_10 = mem_io_portA_output_bits_10; // @[Accumulator.scala 84:13]
  assign io_output_bits_11 = mem_io_portA_output_bits_11; // @[Accumulator.scala 84:13]
  assign io_output_bits_12 = mem_io_portA_output_bits_12; // @[Accumulator.scala 84:13]
  assign io_output_bits_13 = mem_io_portA_output_bits_13; // @[Accumulator.scala 84:13]
  assign io_output_bits_14 = mem_io_portA_output_bits_14; // @[Accumulator.scala 84:13]
  assign io_output_bits_15 = mem_io_portA_output_bits_15; // @[Accumulator.scala 84:13]
  assign io_output_bits_16 = mem_io_portA_output_bits_16; // @[Accumulator.scala 84:13]
  assign io_output_bits_17 = mem_io_portA_output_bits_17; // @[Accumulator.scala 84:13]
  assign io_output_bits_18 = mem_io_portA_output_bits_18; // @[Accumulator.scala 84:13]
  assign io_output_bits_19 = mem_io_portA_output_bits_19; // @[Accumulator.scala 84:13]
  assign io_output_bits_20 = mem_io_portA_output_bits_20; // @[Accumulator.scala 84:13]
  assign io_output_bits_21 = mem_io_portA_output_bits_21; // @[Accumulator.scala 84:13]
  assign io_output_bits_22 = mem_io_portA_output_bits_22; // @[Accumulator.scala 84:13]
  assign io_output_bits_23 = mem_io_portA_output_bits_23; // @[Accumulator.scala 84:13]
  assign io_output_bits_24 = mem_io_portA_output_bits_24; // @[Accumulator.scala 84:13]
  assign io_output_bits_25 = mem_io_portA_output_bits_25; // @[Accumulator.scala 84:13]
  assign io_output_bits_26 = mem_io_portA_output_bits_26; // @[Accumulator.scala 84:13]
  assign io_output_bits_27 = mem_io_portA_output_bits_27; // @[Accumulator.scala 84:13]
  assign io_output_bits_28 = mem_io_portA_output_bits_28; // @[Accumulator.scala 84:13]
  assign io_output_bits_29 = mem_io_portA_output_bits_29; // @[Accumulator.scala 84:13]
  assign io_output_bits_30 = mem_io_portA_output_bits_30; // @[Accumulator.scala 84:13]
  assign io_output_bits_31 = mem_io_portA_output_bits_31; // @[Accumulator.scala 84:13]
  assign io_control_ready = io_control_bits_write ? _GEN_17 : readEnqueuer_io_in_ready; // @[Accumulator.scala 111:28 143:19]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_portA_control_valid = lockPool_io_actor_0_out_valid; // @[Accumulator.scala 66:19]
  assign mem_io_portA_control_bits_write = lockPool_io_actor_0_out_bits_write; // @[Accumulator.scala 66:19]
  assign mem_io_portA_control_bits_address = lockPool_io_actor_0_out_bits_address; // @[Accumulator.scala 66:19]
  assign mem_io_portA_input_valid = portAInputMux_x14_mux_io_out_valid; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_0 = portAInputMux_x14_mux_io_out_bits_0; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_1 = portAInputMux_x14_mux_io_out_bits_1; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_2 = portAInputMux_x14_mux_io_out_bits_2; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_3 = portAInputMux_x14_mux_io_out_bits_3; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_4 = portAInputMux_x14_mux_io_out_bits_4; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_5 = portAInputMux_x14_mux_io_out_bits_5; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_6 = portAInputMux_x14_mux_io_out_bits_6; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_7 = portAInputMux_x14_mux_io_out_bits_7; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_8 = portAInputMux_x14_mux_io_out_bits_8; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_9 = portAInputMux_x14_mux_io_out_bits_9; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_10 = portAInputMux_x14_mux_io_out_bits_10; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_11 = portAInputMux_x14_mux_io_out_bits_11; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_12 = portAInputMux_x14_mux_io_out_bits_12; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_13 = portAInputMux_x14_mux_io_out_bits_13; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_14 = portAInputMux_x14_mux_io_out_bits_14; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_15 = portAInputMux_x14_mux_io_out_bits_15; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_16 = portAInputMux_x14_mux_io_out_bits_16; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_17 = portAInputMux_x14_mux_io_out_bits_17; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_18 = portAInputMux_x14_mux_io_out_bits_18; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_19 = portAInputMux_x14_mux_io_out_bits_19; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_20 = portAInputMux_x14_mux_io_out_bits_20; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_21 = portAInputMux_x14_mux_io_out_bits_21; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_22 = portAInputMux_x14_mux_io_out_bits_22; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_23 = portAInputMux_x14_mux_io_out_bits_23; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_24 = portAInputMux_x14_mux_io_out_bits_24; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_25 = portAInputMux_x14_mux_io_out_bits_25; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_26 = portAInputMux_x14_mux_io_out_bits_26; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_27 = portAInputMux_x14_mux_io_out_bits_27; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_28 = portAInputMux_x14_mux_io_out_bits_28; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_29 = portAInputMux_x14_mux_io_out_bits_29; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_30 = portAInputMux_x14_mux_io_out_bits_30; // @[Mux.scala 81:9]
  assign mem_io_portA_input_bits_31 = portAInputMux_x14_mux_io_out_bits_31; // @[Mux.scala 81:9]
  assign mem_io_portA_output_ready = io_output_ready; // @[Accumulator.scala 84:13]
  assign mem_io_portB_control_valid = lockPool_io_actor_1_out_valid; // @[Accumulator.scala 67:19]
  assign mem_io_portB_control_bits_address = lockPool_io_actor_1_out_bits_address; // @[Accumulator.scala 67:19]
  assign mem_io_portB_output_ready = adder_io_right_ready; // @[Accumulator.scala 86:18]
  assign mem_io_tracepoint = io_tracepoint; // @[Accumulator.scala 74:21]
  assign mem_io_programCounter = io_programCounter; // @[Accumulator.scala 73:25]
  assign adder_io_left_valid = inputDemuxModule_io_out_1_valid; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_0 = inputDemuxModule_io_out_1_bits_0; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_1 = inputDemuxModule_io_out_1_bits_1; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_2 = inputDemuxModule_io_out_1_bits_2; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_3 = inputDemuxModule_io_out_1_bits_3; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_4 = inputDemuxModule_io_out_1_bits_4; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_5 = inputDemuxModule_io_out_1_bits_5; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_6 = inputDemuxModule_io_out_1_bits_6; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_7 = inputDemuxModule_io_out_1_bits_7; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_8 = inputDemuxModule_io_out_1_bits_8; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_9 = inputDemuxModule_io_out_1_bits_9; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_10 = inputDemuxModule_io_out_1_bits_10; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_11 = inputDemuxModule_io_out_1_bits_11; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_12 = inputDemuxModule_io_out_1_bits_12; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_13 = inputDemuxModule_io_out_1_bits_13; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_14 = inputDemuxModule_io_out_1_bits_14; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_15 = inputDemuxModule_io_out_1_bits_15; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_16 = inputDemuxModule_io_out_1_bits_16; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_17 = inputDemuxModule_io_out_1_bits_17; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_18 = inputDemuxModule_io_out_1_bits_18; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_19 = inputDemuxModule_io_out_1_bits_19; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_20 = inputDemuxModule_io_out_1_bits_20; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_21 = inputDemuxModule_io_out_1_bits_21; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_22 = inputDemuxModule_io_out_1_bits_22; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_23 = inputDemuxModule_io_out_1_bits_23; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_24 = inputDemuxModule_io_out_1_bits_24; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_25 = inputDemuxModule_io_out_1_bits_25; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_26 = inputDemuxModule_io_out_1_bits_26; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_27 = inputDemuxModule_io_out_1_bits_27; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_28 = inputDemuxModule_io_out_1_bits_28; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_29 = inputDemuxModule_io_out_1_bits_29; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_30 = inputDemuxModule_io_out_1_bits_30; // @[Accumulator.scala 94:17]
  assign adder_io_left_bits_31 = inputDemuxModule_io_out_1_bits_31; // @[Accumulator.scala 94:17]
  assign adder_io_right_valid = mem_io_portB_output_valid; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_0 = mem_io_portB_output_bits_0; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_1 = mem_io_portB_output_bits_1; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_2 = mem_io_portB_output_bits_2; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_3 = mem_io_portB_output_bits_3; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_4 = mem_io_portB_output_bits_4; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_5 = mem_io_portB_output_bits_5; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_6 = mem_io_portB_output_bits_6; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_7 = mem_io_portB_output_bits_7; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_8 = mem_io_portB_output_bits_8; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_9 = mem_io_portB_output_bits_9; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_10 = mem_io_portB_output_bits_10; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_11 = mem_io_portB_output_bits_11; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_12 = mem_io_portB_output_bits_12; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_13 = mem_io_portB_output_bits_13; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_14 = mem_io_portB_output_bits_14; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_15 = mem_io_portB_output_bits_15; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_16 = mem_io_portB_output_bits_16; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_17 = mem_io_portB_output_bits_17; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_18 = mem_io_portB_output_bits_18; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_19 = mem_io_portB_output_bits_19; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_20 = mem_io_portB_output_bits_20; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_21 = mem_io_portB_output_bits_21; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_22 = mem_io_portB_output_bits_22; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_23 = mem_io_portB_output_bits_23; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_24 = mem_io_portB_output_bits_24; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_25 = mem_io_portB_output_bits_25; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_26 = mem_io_portB_output_bits_26; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_27 = mem_io_portB_output_bits_27; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_28 = mem_io_portB_output_bits_28; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_29 = mem_io_portB_output_bits_29; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_30 = mem_io_portB_output_bits_30; // @[Accumulator.scala 86:18]
  assign adder_io_right_bits_31 = mem_io_portB_output_bits_31; // @[Accumulator.scala 86:18]
  assign adder_io_output_ready = portAInputMux_x14_mux_io_in_1_ready; // @[Mux.scala 80:18]
  assign lockPool_clock = clock;
  assign lockPool_reset = reset;
  assign lockPool_io_actor_0_in_valid = portAControl_io_deq_valid; // @[Mem.scala 23:7]
  assign lockPool_io_actor_0_in_bits_write = portAControl_io_deq_bits_write; // @[Mem.scala 23:7]
  assign lockPool_io_actor_0_in_bits_address = portAControl_io_deq_bits_address; // @[Mem.scala 23:7]
  assign lockPool_io_actor_0_in_bits_size = portAControl_io_deq_bits_size; // @[Mem.scala 23:7]
  assign lockPool_io_actor_0_out_ready = mem_io_portA_control_ready; // @[Accumulator.scala 66:19]
  assign lockPool_io_actor_1_in_valid = io_control_bits_write & _GEN_7; // @[Accumulator.scala 111:28 package.scala 405:15]
  assign lockPool_io_actor_1_in_bits_address = io_control_bits_write ? _GEN_9 : 12'h0; // @[Accumulator.scala 111:28 package.scala 404:14]
  assign lockPool_io_actor_1_out_ready = mem_io_portB_control_ready; // @[Accumulator.scala 67:19]
  assign lockPool_io_lock_valid = io_control_bits_write & _GEN_23; // @[Accumulator.scala 111:28 Decoupled.scala 72:20]
  assign lockPool_io_lock_bits_cond_address = io_control_bits_address; // @[MemControl.scala 67:17 68:15]
  assign portAControl_clock = clock;
  assign portAControl_reset = reset;
  assign portAControl_io_enq_valid = io_control_bits_write ? _GEN_2 : io_control_ready_portAControl_io_enq_w_2_valid; // @[Accumulator.scala 111:28 MultiEnqueue.scala 61:10]
  assign portAControl_io_enq_bits_write = io_control_bits_write; // @[Accumulator.scala 111:28 MultiEnqueue.scala 61:10]
  assign portAControl_io_enq_bits_address = io_control_bits_address; // @[Accumulator.scala 111:28 MultiEnqueue.scala 61:10]
  assign portAControl_io_deq_ready = lockPool_io_actor_0_in_ready; // @[Mem.scala 23:7]
  assign inputDemuxModule_io_in_valid = io_input_valid; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_0 = io_input_bits_0; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_1 = io_input_bits_1; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_2 = io_input_bits_2; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_3 = io_input_bits_3; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_4 = io_input_bits_4; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_5 = io_input_bits_5; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_6 = io_input_bits_6; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_7 = io_input_bits_7; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_8 = io_input_bits_8; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_9 = io_input_bits_9; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_10 = io_input_bits_10; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_11 = io_input_bits_11; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_12 = io_input_bits_12; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_13 = io_input_bits_13; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_14 = io_input_bits_14; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_15 = io_input_bits_15; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_16 = io_input_bits_16; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_17 = io_input_bits_17; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_18 = io_input_bits_18; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_19 = io_input_bits_19; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_20 = io_input_bits_20; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_21 = io_input_bits_21; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_22 = io_input_bits_22; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_23 = io_input_bits_23; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_24 = io_input_bits_24; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_25 = io_input_bits_25; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_26 = io_input_bits_26; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_27 = io_input_bits_27; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_28 = io_input_bits_28; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_29 = io_input_bits_29; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_30 = io_input_bits_30; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_in_bits_31 = io_input_bits_31; // @[Accumulator.scala 93:26]
  assign inputDemuxModule_io_sel_valid = inputDemux_io_deq_valid; // @[Mem.scala 23:7]
  assign inputDemuxModule_io_sel_bits = inputDemux_io_deq_bits; // @[Mem.scala 23:7]
  assign inputDemuxModule_io_out_0_ready = portAInputMux_x14_mux_io_in_0_ready; // @[Mux.scala 79:18]
  assign inputDemuxModule_io_out_1_ready = adder_io_left_ready; // @[Accumulator.scala 94:17]
  assign inputDemux_clock = clock;
  assign inputDemux_reset = reset;
  assign inputDemux_io_enq_valid = io_control_bits_write & _GEN_12; // @[Accumulator.scala 111:28 Decoupled.scala 72:20]
  assign inputDemux_io_enq_bits = io_control_bits_accumulate; // @[Accumulator.scala 112:35 MultiEnqueue.scala 152:10 153:10]
  assign inputDemux_io_deq_ready = inputDemuxModule_io_sel_ready; // @[Mem.scala 23:7]
  assign portAInputMux_x14_mux_io_in_0_valid = inputDemuxModule_io_out_0_valid; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_0 = inputDemuxModule_io_out_0_bits_0; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_1 = inputDemuxModule_io_out_0_bits_1; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_2 = inputDemuxModule_io_out_0_bits_2; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_3 = inputDemuxModule_io_out_0_bits_3; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_4 = inputDemuxModule_io_out_0_bits_4; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_5 = inputDemuxModule_io_out_0_bits_5; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_6 = inputDemuxModule_io_out_0_bits_6; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_7 = inputDemuxModule_io_out_0_bits_7; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_8 = inputDemuxModule_io_out_0_bits_8; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_9 = inputDemuxModule_io_out_0_bits_9; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_10 = inputDemuxModule_io_out_0_bits_10; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_11 = inputDemuxModule_io_out_0_bits_11; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_12 = inputDemuxModule_io_out_0_bits_12; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_13 = inputDemuxModule_io_out_0_bits_13; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_14 = inputDemuxModule_io_out_0_bits_14; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_15 = inputDemuxModule_io_out_0_bits_15; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_16 = inputDemuxModule_io_out_0_bits_16; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_17 = inputDemuxModule_io_out_0_bits_17; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_18 = inputDemuxModule_io_out_0_bits_18; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_19 = inputDemuxModule_io_out_0_bits_19; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_20 = inputDemuxModule_io_out_0_bits_20; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_21 = inputDemuxModule_io_out_0_bits_21; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_22 = inputDemuxModule_io_out_0_bits_22; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_23 = inputDemuxModule_io_out_0_bits_23; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_24 = inputDemuxModule_io_out_0_bits_24; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_25 = inputDemuxModule_io_out_0_bits_25; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_26 = inputDemuxModule_io_out_0_bits_26; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_27 = inputDemuxModule_io_out_0_bits_27; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_28 = inputDemuxModule_io_out_0_bits_28; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_29 = inputDemuxModule_io_out_0_bits_29; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_30 = inputDemuxModule_io_out_0_bits_30; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_0_bits_31 = inputDemuxModule_io_out_0_bits_31; // @[Mux.scala 79:18]
  assign portAInputMux_x14_mux_io_in_1_valid = adder_io_output_valid; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_0 = adder_io_output_bits_0; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_1 = adder_io_output_bits_1; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_2 = adder_io_output_bits_2; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_3 = adder_io_output_bits_3; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_4 = adder_io_output_bits_4; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_5 = adder_io_output_bits_5; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_6 = adder_io_output_bits_6; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_7 = adder_io_output_bits_7; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_8 = adder_io_output_bits_8; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_9 = adder_io_output_bits_9; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_10 = adder_io_output_bits_10; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_11 = adder_io_output_bits_11; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_12 = adder_io_output_bits_12; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_13 = adder_io_output_bits_13; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_14 = adder_io_output_bits_14; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_15 = adder_io_output_bits_15; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_16 = adder_io_output_bits_16; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_17 = adder_io_output_bits_17; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_18 = adder_io_output_bits_18; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_19 = adder_io_output_bits_19; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_20 = adder_io_output_bits_20; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_21 = adder_io_output_bits_21; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_22 = adder_io_output_bits_22; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_23 = adder_io_output_bits_23; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_24 = adder_io_output_bits_24; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_25 = adder_io_output_bits_25; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_26 = adder_io_output_bits_26; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_27 = adder_io_output_bits_27; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_28 = adder_io_output_bits_28; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_29 = adder_io_output_bits_29; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_30 = adder_io_output_bits_30; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_in_1_bits_31 = adder_io_output_bits_31; // @[Mux.scala 80:18]
  assign portAInputMux_x14_mux_io_sel_valid = portAInputMux_io_deq_valid; // @[Mem.scala 23:7]
  assign portAInputMux_x14_mux_io_sel_bits = portAInputMux_io_deq_bits; // @[Mem.scala 23:7]
  assign portAInputMux_x14_mux_io_out_ready = mem_io_portA_input_ready; // @[Mux.scala 81:9]
  assign portAInputMux_clock = clock;
  assign portAInputMux_reset = reset;
  assign portAInputMux_io_enq_valid = io_control_bits_write & _GEN_15; // @[Accumulator.scala 111:28 Decoupled.scala 72:20]
  assign portAInputMux_io_enq_bits = io_control_bits_accumulate; // @[Accumulator.scala 112:35 MultiEnqueue.scala 153:10 154:10]
  assign portAInputMux_io_deq_ready = portAInputMux_x14_mux_io_sel_ready; // @[Mem.scala 23:7]
  assign writeEnqueuer_clock = clock;
  assign writeEnqueuer_reset = reset;
  assign writeEnqueuer_io_in_valid = io_control_bits_write & _GEN_18; // @[Accumulator.scala 111:28 MultiEnqueue.scala 40:17]
  assign writeEnqueuer_io_out_0_ready = io_control_bits_write & _GEN_19; // @[Accumulator.scala 111:28 MultiEnqueue.scala 42:18]
  assign writeEnqueuer_io_out_1_ready = io_control_bits_write & _GEN_20; // @[Accumulator.scala 111:28 MultiEnqueue.scala 42:18]
  assign writeEnqueuer_io_out_2_ready = io_control_bits_write & _GEN_21; // @[Accumulator.scala 111:28 MultiEnqueue.scala 42:18]
  assign writeEnqueuer_io_out_3_ready = io_control_bits_write & _GEN_22; // @[Accumulator.scala 111:28 MultiEnqueue.scala 42:18]
  assign readEnqueuer_clock = clock;
  assign readEnqueuer_reset = reset;
  assign readEnqueuer_io_in_valid = io_control_bits_write ? 1'h0 : io_control_valid; // @[Accumulator.scala 111:28 MultiEnqueue.scala 40:17 60:17]
  assign readEnqueuer_io_out_0_ready = io_control_bits_write ? 1'h0 : io_control_ready_portAControl_io_enq_w_ready; // @[Accumulator.scala 111:28 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  assign accEnqueuer_clock = clock;
  assign accEnqueuer_reset = reset;
  assign accEnqueuer_io_in_valid = io_control_bits_write & _GEN_0; // @[Accumulator.scala 111:28 MultiEnqueue.scala 40:17]
  assign accEnqueuer_io_out_0_ready = io_control_bits_write & _GEN_1; // @[Accumulator.scala 111:28 MultiEnqueue.scala 42:18]
  assign accEnqueuer_io_out_1_ready = io_control_bits_write & _GEN_6; // @[Accumulator.scala 111:28 MultiEnqueue.scala 42:18]
  assign accEnqueuer_io_out_2_ready = io_control_bits_write & _GEN_11; // @[Accumulator.scala 111:28 MultiEnqueue.scala 42:18]
  assign accEnqueuer_io_out_3_ready = io_control_bits_write & _GEN_14; // @[Accumulator.scala 111:28 MultiEnqueue.scala 42:18]
endmodule
module Queue_17(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_0,
  input  [15:0] io_enq_bits_1,
  input  [15:0] io_enq_bits_2,
  input  [15:0] io_enq_bits_3,
  input  [15:0] io_enq_bits_4,
  input  [15:0] io_enq_bits_5,
  input  [15:0] io_enq_bits_6,
  input  [15:0] io_enq_bits_7,
  input  [15:0] io_enq_bits_8,
  input  [15:0] io_enq_bits_9,
  input  [15:0] io_enq_bits_10,
  input  [15:0] io_enq_bits_11,
  input  [15:0] io_enq_bits_12,
  input  [15:0] io_enq_bits_13,
  input  [15:0] io_enq_bits_14,
  input  [15:0] io_enq_bits_15,
  input  [15:0] io_enq_bits_16,
  input  [15:0] io_enq_bits_17,
  input  [15:0] io_enq_bits_18,
  input  [15:0] io_enq_bits_19,
  input  [15:0] io_enq_bits_20,
  input  [15:0] io_enq_bits_21,
  input  [15:0] io_enq_bits_22,
  input  [15:0] io_enq_bits_23,
  input  [15:0] io_enq_bits_24,
  input  [15:0] io_enq_bits_25,
  input  [15:0] io_enq_bits_26,
  input  [15:0] io_enq_bits_27,
  input  [15:0] io_enq_bits_28,
  input  [15:0] io_enq_bits_29,
  input  [15:0] io_enq_bits_30,
  input  [15:0] io_enq_bits_31,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_0,
  output [15:0] io_deq_bits_1,
  output [15:0] io_deq_bits_2,
  output [15:0] io_deq_bits_3,
  output [15:0] io_deq_bits_4,
  output [15:0] io_deq_bits_5,
  output [15:0] io_deq_bits_6,
  output [15:0] io_deq_bits_7,
  output [15:0] io_deq_bits_8,
  output [15:0] io_deq_bits_9,
  output [15:0] io_deq_bits_10,
  output [15:0] io_deq_bits_11,
  output [15:0] io_deq_bits_12,
  output [15:0] io_deq_bits_13,
  output [15:0] io_deq_bits_14,
  output [15:0] io_deq_bits_15,
  output [15:0] io_deq_bits_16,
  output [15:0] io_deq_bits_17,
  output [15:0] io_deq_bits_18,
  output [15:0] io_deq_bits_19,
  output [15:0] io_deq_bits_20,
  output [15:0] io_deq_bits_21,
  output [15:0] io_deq_bits_22,
  output [15:0] io_deq_bits_23,
  output [15:0] io_deq_bits_24,
  output [15:0] io_deq_bits_25,
  output [15:0] io_deq_bits_26,
  output [15:0] io_deq_bits_27,
  output [15:0] io_deq_bits_28,
  output [15:0] io_deq_bits_29,
  output [15:0] io_deq_bits_30,
  output [15:0] io_deq_bits_31
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ram_0 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_1 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_2 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_3 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_4 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_5 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_6 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_7 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_8 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_8_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_8_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_8_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_8_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_8_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_8_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_8_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_9 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_9_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_9_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_9_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_9_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_9_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_9_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_9_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_10 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_10_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_10_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_10_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_10_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_10_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_10_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_10_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_11 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_11_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_11_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_11_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_11_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_11_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_11_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_11_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_12 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_12_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_12_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_12_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_12_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_12_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_12_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_12_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_13 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_13_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_13_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_13_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_13_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_13_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_13_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_13_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_14 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_14_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_14_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_14_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_14_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_14_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_14_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_14_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_15 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_15_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_15_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_15_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_15_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_15_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_15_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_15_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_16 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_16_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_16_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_16_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_16_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_16_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_16_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_16_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_17 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_17_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_17_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_17_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_17_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_17_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_17_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_17_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_18 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_18_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_18_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_18_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_18_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_18_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_18_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_18_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_19 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_19_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_19_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_19_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_19_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_19_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_19_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_19_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_20 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_20_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_20_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_20_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_20_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_20_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_20_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_20_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_21 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_21_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_21_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_21_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_21_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_21_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_21_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_21_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_22 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_22_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_22_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_22_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_22_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_22_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_22_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_22_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_23 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_23_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_23_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_23_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_23_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_23_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_23_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_23_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_24 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_24_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_24_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_24_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_24_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_24_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_24_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_24_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_25 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_25_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_25_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_25_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_25_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_25_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_25_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_25_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_26 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_26_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_26_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_26_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_26_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_26_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_26_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_26_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_27 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_27_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_27_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_27_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_27_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_27_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_27_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_27_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_28 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_28_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_28_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_28_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_28_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_28_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_28_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_28_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_29 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_29_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_29_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_29_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_29_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_29_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_29_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_29_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_30 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_30_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_30_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_30_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_30_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_30_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_30_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_30_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_31 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_31_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_31_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_31_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_31_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_31_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_31_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_31_MPORT_en; // @[Decoupled.scala 259:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_43 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_43 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_0_io_deq_bits_MPORT_data = ram_0[ram_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_0_MPORT_data = io_enq_bits_0;
  assign ram_0_MPORT_addr = enq_ptr_value;
  assign ram_0_MPORT_mask = 1'h1;
  assign ram_0_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_1_io_deq_bits_MPORT_data = ram_1[ram_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_1_MPORT_data = io_enq_bits_1;
  assign ram_1_MPORT_addr = enq_ptr_value;
  assign ram_1_MPORT_mask = 1'h1;
  assign ram_1_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_2_io_deq_bits_MPORT_data = ram_2[ram_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_2_MPORT_data = io_enq_bits_2;
  assign ram_2_MPORT_addr = enq_ptr_value;
  assign ram_2_MPORT_mask = 1'h1;
  assign ram_2_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_3_io_deq_bits_MPORT_data = ram_3[ram_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_3_MPORT_data = io_enq_bits_3;
  assign ram_3_MPORT_addr = enq_ptr_value;
  assign ram_3_MPORT_mask = 1'h1;
  assign ram_3_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_4_io_deq_bits_MPORT_data = ram_4[ram_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_4_MPORT_data = io_enq_bits_4;
  assign ram_4_MPORT_addr = enq_ptr_value;
  assign ram_4_MPORT_mask = 1'h1;
  assign ram_4_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_5_io_deq_bits_MPORT_data = ram_5[ram_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_5_MPORT_data = io_enq_bits_5;
  assign ram_5_MPORT_addr = enq_ptr_value;
  assign ram_5_MPORT_mask = 1'h1;
  assign ram_5_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_6_io_deq_bits_MPORT_data = ram_6[ram_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_6_MPORT_data = io_enq_bits_6;
  assign ram_6_MPORT_addr = enq_ptr_value;
  assign ram_6_MPORT_mask = 1'h1;
  assign ram_6_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_7_io_deq_bits_MPORT_data = ram_7[ram_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_7_MPORT_data = io_enq_bits_7;
  assign ram_7_MPORT_addr = enq_ptr_value;
  assign ram_7_MPORT_mask = 1'h1;
  assign ram_7_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_8_io_deq_bits_MPORT_en = 1'h1;
  assign ram_8_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_8_io_deq_bits_MPORT_data = ram_8[ram_8_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_8_MPORT_data = io_enq_bits_8;
  assign ram_8_MPORT_addr = enq_ptr_value;
  assign ram_8_MPORT_mask = 1'h1;
  assign ram_8_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_9_io_deq_bits_MPORT_en = 1'h1;
  assign ram_9_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_9_io_deq_bits_MPORT_data = ram_9[ram_9_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_9_MPORT_data = io_enq_bits_9;
  assign ram_9_MPORT_addr = enq_ptr_value;
  assign ram_9_MPORT_mask = 1'h1;
  assign ram_9_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_10_io_deq_bits_MPORT_en = 1'h1;
  assign ram_10_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_10_io_deq_bits_MPORT_data = ram_10[ram_10_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_10_MPORT_data = io_enq_bits_10;
  assign ram_10_MPORT_addr = enq_ptr_value;
  assign ram_10_MPORT_mask = 1'h1;
  assign ram_10_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_11_io_deq_bits_MPORT_en = 1'h1;
  assign ram_11_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_11_io_deq_bits_MPORT_data = ram_11[ram_11_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_11_MPORT_data = io_enq_bits_11;
  assign ram_11_MPORT_addr = enq_ptr_value;
  assign ram_11_MPORT_mask = 1'h1;
  assign ram_11_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_12_io_deq_bits_MPORT_en = 1'h1;
  assign ram_12_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_12_io_deq_bits_MPORT_data = ram_12[ram_12_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_12_MPORT_data = io_enq_bits_12;
  assign ram_12_MPORT_addr = enq_ptr_value;
  assign ram_12_MPORT_mask = 1'h1;
  assign ram_12_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_13_io_deq_bits_MPORT_en = 1'h1;
  assign ram_13_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_13_io_deq_bits_MPORT_data = ram_13[ram_13_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_13_MPORT_data = io_enq_bits_13;
  assign ram_13_MPORT_addr = enq_ptr_value;
  assign ram_13_MPORT_mask = 1'h1;
  assign ram_13_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_14_io_deq_bits_MPORT_en = 1'h1;
  assign ram_14_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_14_io_deq_bits_MPORT_data = ram_14[ram_14_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_14_MPORT_data = io_enq_bits_14;
  assign ram_14_MPORT_addr = enq_ptr_value;
  assign ram_14_MPORT_mask = 1'h1;
  assign ram_14_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_15_io_deq_bits_MPORT_en = 1'h1;
  assign ram_15_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_15_io_deq_bits_MPORT_data = ram_15[ram_15_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_15_MPORT_data = io_enq_bits_15;
  assign ram_15_MPORT_addr = enq_ptr_value;
  assign ram_15_MPORT_mask = 1'h1;
  assign ram_15_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_16_io_deq_bits_MPORT_en = 1'h1;
  assign ram_16_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_16_io_deq_bits_MPORT_data = ram_16[ram_16_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_16_MPORT_data = io_enq_bits_16;
  assign ram_16_MPORT_addr = enq_ptr_value;
  assign ram_16_MPORT_mask = 1'h1;
  assign ram_16_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_17_io_deq_bits_MPORT_en = 1'h1;
  assign ram_17_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_17_io_deq_bits_MPORT_data = ram_17[ram_17_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_17_MPORT_data = io_enq_bits_17;
  assign ram_17_MPORT_addr = enq_ptr_value;
  assign ram_17_MPORT_mask = 1'h1;
  assign ram_17_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_18_io_deq_bits_MPORT_en = 1'h1;
  assign ram_18_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_18_io_deq_bits_MPORT_data = ram_18[ram_18_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_18_MPORT_data = io_enq_bits_18;
  assign ram_18_MPORT_addr = enq_ptr_value;
  assign ram_18_MPORT_mask = 1'h1;
  assign ram_18_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_19_io_deq_bits_MPORT_en = 1'h1;
  assign ram_19_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_19_io_deq_bits_MPORT_data = ram_19[ram_19_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_19_MPORT_data = io_enq_bits_19;
  assign ram_19_MPORT_addr = enq_ptr_value;
  assign ram_19_MPORT_mask = 1'h1;
  assign ram_19_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_20_io_deq_bits_MPORT_en = 1'h1;
  assign ram_20_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_20_io_deq_bits_MPORT_data = ram_20[ram_20_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_20_MPORT_data = io_enq_bits_20;
  assign ram_20_MPORT_addr = enq_ptr_value;
  assign ram_20_MPORT_mask = 1'h1;
  assign ram_20_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_21_io_deq_bits_MPORT_en = 1'h1;
  assign ram_21_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_21_io_deq_bits_MPORT_data = ram_21[ram_21_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_21_MPORT_data = io_enq_bits_21;
  assign ram_21_MPORT_addr = enq_ptr_value;
  assign ram_21_MPORT_mask = 1'h1;
  assign ram_21_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_22_io_deq_bits_MPORT_en = 1'h1;
  assign ram_22_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_22_io_deq_bits_MPORT_data = ram_22[ram_22_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_22_MPORT_data = io_enq_bits_22;
  assign ram_22_MPORT_addr = enq_ptr_value;
  assign ram_22_MPORT_mask = 1'h1;
  assign ram_22_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_23_io_deq_bits_MPORT_en = 1'h1;
  assign ram_23_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_23_io_deq_bits_MPORT_data = ram_23[ram_23_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_23_MPORT_data = io_enq_bits_23;
  assign ram_23_MPORT_addr = enq_ptr_value;
  assign ram_23_MPORT_mask = 1'h1;
  assign ram_23_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_24_io_deq_bits_MPORT_en = 1'h1;
  assign ram_24_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_24_io_deq_bits_MPORT_data = ram_24[ram_24_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_24_MPORT_data = io_enq_bits_24;
  assign ram_24_MPORT_addr = enq_ptr_value;
  assign ram_24_MPORT_mask = 1'h1;
  assign ram_24_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_25_io_deq_bits_MPORT_en = 1'h1;
  assign ram_25_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_25_io_deq_bits_MPORT_data = ram_25[ram_25_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_25_MPORT_data = io_enq_bits_25;
  assign ram_25_MPORT_addr = enq_ptr_value;
  assign ram_25_MPORT_mask = 1'h1;
  assign ram_25_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_26_io_deq_bits_MPORT_en = 1'h1;
  assign ram_26_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_26_io_deq_bits_MPORT_data = ram_26[ram_26_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_26_MPORT_data = io_enq_bits_26;
  assign ram_26_MPORT_addr = enq_ptr_value;
  assign ram_26_MPORT_mask = 1'h1;
  assign ram_26_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_27_io_deq_bits_MPORT_en = 1'h1;
  assign ram_27_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_27_io_deq_bits_MPORT_data = ram_27[ram_27_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_27_MPORT_data = io_enq_bits_27;
  assign ram_27_MPORT_addr = enq_ptr_value;
  assign ram_27_MPORT_mask = 1'h1;
  assign ram_27_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_28_io_deq_bits_MPORT_en = 1'h1;
  assign ram_28_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_28_io_deq_bits_MPORT_data = ram_28[ram_28_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_28_MPORT_data = io_enq_bits_28;
  assign ram_28_MPORT_addr = enq_ptr_value;
  assign ram_28_MPORT_mask = 1'h1;
  assign ram_28_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_29_io_deq_bits_MPORT_en = 1'h1;
  assign ram_29_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_29_io_deq_bits_MPORT_data = ram_29[ram_29_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_29_MPORT_data = io_enq_bits_29;
  assign ram_29_MPORT_addr = enq_ptr_value;
  assign ram_29_MPORT_mask = 1'h1;
  assign ram_29_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_30_io_deq_bits_MPORT_en = 1'h1;
  assign ram_30_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_30_io_deq_bits_MPORT_data = ram_30[ram_30_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_30_MPORT_data = io_enq_bits_30;
  assign ram_30_MPORT_addr = enq_ptr_value;
  assign ram_30_MPORT_mask = 1'h1;
  assign ram_30_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign ram_31_io_deq_bits_MPORT_en = 1'h1;
  assign ram_31_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_31_io_deq_bits_MPORT_data = ram_31[ram_31_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_31_MPORT_data = io_enq_bits_31;
  assign ram_31_MPORT_addr = enq_ptr_value;
  assign ram_31_MPORT_mask = 1'h1;
  assign ram_31_MPORT_en = empty ? _GEN_43 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_0 = empty ? $signed(io_enq_bits_0) : $signed(ram_0_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_1 = empty ? $signed(io_enq_bits_1) : $signed(ram_1_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_2 = empty ? $signed(io_enq_bits_2) : $signed(ram_2_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_3 = empty ? $signed(io_enq_bits_3) : $signed(ram_3_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_4 = empty ? $signed(io_enq_bits_4) : $signed(ram_4_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_5 = empty ? $signed(io_enq_bits_5) : $signed(ram_5_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_6 = empty ? $signed(io_enq_bits_6) : $signed(ram_6_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_7 = empty ? $signed(io_enq_bits_7) : $signed(ram_7_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_8 = empty ? $signed(io_enq_bits_8) : $signed(ram_8_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_9 = empty ? $signed(io_enq_bits_9) : $signed(ram_9_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_10 = empty ? $signed(io_enq_bits_10) : $signed(ram_10_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_11 = empty ? $signed(io_enq_bits_11) : $signed(ram_11_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_12 = empty ? $signed(io_enq_bits_12) : $signed(ram_12_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_13 = empty ? $signed(io_enq_bits_13) : $signed(ram_13_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_14 = empty ? $signed(io_enq_bits_14) : $signed(ram_14_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_15 = empty ? $signed(io_enq_bits_15) : $signed(ram_15_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_16 = empty ? $signed(io_enq_bits_16) : $signed(ram_16_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_17 = empty ? $signed(io_enq_bits_17) : $signed(ram_17_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_18 = empty ? $signed(io_enq_bits_18) : $signed(ram_18_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_19 = empty ? $signed(io_enq_bits_19) : $signed(ram_19_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_20 = empty ? $signed(io_enq_bits_20) : $signed(ram_20_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_21 = empty ? $signed(io_enq_bits_21) : $signed(ram_21_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_22 = empty ? $signed(io_enq_bits_22) : $signed(ram_22_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_23 = empty ? $signed(io_enq_bits_23) : $signed(ram_23_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_24 = empty ? $signed(io_enq_bits_24) : $signed(ram_24_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_25 = empty ? $signed(io_enq_bits_25) : $signed(ram_25_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_26 = empty ? $signed(io_enq_bits_26) : $signed(ram_26_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_27 = empty ? $signed(io_enq_bits_27) : $signed(ram_27_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_28 = empty ? $signed(io_enq_bits_28) : $signed(ram_28_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_29 = empty ? $signed(io_enq_bits_29) : $signed(ram_29_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_30 = empty ? $signed(io_enq_bits_30) : $signed(ram_30_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_31 = empty ? $signed(io_enq_bits_31) : $signed(ram_31_io_deq_bits_MPORT_data); // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_0_MPORT_en & ram_0_MPORT_mask) begin
      ram_0[ram_0_MPORT_addr] <= ram_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_1_MPORT_en & ram_1_MPORT_mask) begin
      ram_1[ram_1_MPORT_addr] <= ram_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_2_MPORT_en & ram_2_MPORT_mask) begin
      ram_2[ram_2_MPORT_addr] <= ram_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_3_MPORT_en & ram_3_MPORT_mask) begin
      ram_3[ram_3_MPORT_addr] <= ram_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_4_MPORT_en & ram_4_MPORT_mask) begin
      ram_4[ram_4_MPORT_addr] <= ram_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_5_MPORT_en & ram_5_MPORT_mask) begin
      ram_5[ram_5_MPORT_addr] <= ram_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_6_MPORT_en & ram_6_MPORT_mask) begin
      ram_6[ram_6_MPORT_addr] <= ram_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_7_MPORT_en & ram_7_MPORT_mask) begin
      ram_7[ram_7_MPORT_addr] <= ram_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_8_MPORT_en & ram_8_MPORT_mask) begin
      ram_8[ram_8_MPORT_addr] <= ram_8_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_9_MPORT_en & ram_9_MPORT_mask) begin
      ram_9[ram_9_MPORT_addr] <= ram_9_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_10_MPORT_en & ram_10_MPORT_mask) begin
      ram_10[ram_10_MPORT_addr] <= ram_10_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_11_MPORT_en & ram_11_MPORT_mask) begin
      ram_11[ram_11_MPORT_addr] <= ram_11_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_12_MPORT_en & ram_12_MPORT_mask) begin
      ram_12[ram_12_MPORT_addr] <= ram_12_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_13_MPORT_en & ram_13_MPORT_mask) begin
      ram_13[ram_13_MPORT_addr] <= ram_13_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_14_MPORT_en & ram_14_MPORT_mask) begin
      ram_14[ram_14_MPORT_addr] <= ram_14_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_15_MPORT_en & ram_15_MPORT_mask) begin
      ram_15[ram_15_MPORT_addr] <= ram_15_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_16_MPORT_en & ram_16_MPORT_mask) begin
      ram_16[ram_16_MPORT_addr] <= ram_16_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_17_MPORT_en & ram_17_MPORT_mask) begin
      ram_17[ram_17_MPORT_addr] <= ram_17_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_18_MPORT_en & ram_18_MPORT_mask) begin
      ram_18[ram_18_MPORT_addr] <= ram_18_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_19_MPORT_en & ram_19_MPORT_mask) begin
      ram_19[ram_19_MPORT_addr] <= ram_19_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_20_MPORT_en & ram_20_MPORT_mask) begin
      ram_20[ram_20_MPORT_addr] <= ram_20_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_21_MPORT_en & ram_21_MPORT_mask) begin
      ram_21[ram_21_MPORT_addr] <= ram_21_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_22_MPORT_en & ram_22_MPORT_mask) begin
      ram_22[ram_22_MPORT_addr] <= ram_22_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_23_MPORT_en & ram_23_MPORT_mask) begin
      ram_23[ram_23_MPORT_addr] <= ram_23_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_24_MPORT_en & ram_24_MPORT_mask) begin
      ram_24[ram_24_MPORT_addr] <= ram_24_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_25_MPORT_en & ram_25_MPORT_mask) begin
      ram_25[ram_25_MPORT_addr] <= ram_25_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_26_MPORT_en & ram_26_MPORT_mask) begin
      ram_26[ram_26_MPORT_addr] <= ram_26_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_27_MPORT_en & ram_27_MPORT_mask) begin
      ram_27[ram_27_MPORT_addr] <= ram_27_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_28_MPORT_en & ram_28_MPORT_mask) begin
      ram_28[ram_28_MPORT_addr] <= ram_28_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_29_MPORT_en & ram_29_MPORT_mask) begin
      ram_29[ram_29_MPORT_addr] <= ram_29_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_30_MPORT_en & ram_30_MPORT_mask) begin
      ram_30[ram_30_MPORT_addr] <= ram_30_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_31_MPORT_en & ram_31_MPORT_mask) begin
      ram_31[ram_31_MPORT_addr] <= ram_31_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_0[initvar] = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_1[initvar] = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_2[initvar] = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_3[initvar] = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_4[initvar] = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_5[initvar] = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_6[initvar] = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_7[initvar] = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_8[initvar] = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_9[initvar] = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_10[initvar] = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_11[initvar] = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_12[initvar] = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_13[initvar] = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_14[initvar] = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_15[initvar] = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_16[initvar] = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_17[initvar] = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_18[initvar] = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_19[initvar] = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_20[initvar] = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_21[initvar] = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_22[initvar] = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_23[initvar] = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_24[initvar] = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_25[initvar] = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_26[initvar] = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_27[initvar] = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_28[initvar] = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_29[initvar] = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_30[initvar] = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_31[initvar] = _RAND_31[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  enq_ptr_value = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  deq_ptr_value = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  maybe_full = _RAND_34[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [3:0]  io_op,
  input  [15:0] io_input,
  input         io_sourceLeft,
  input         io_sourceRight,
  input         io_dest,
  output [15:0] io_output
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] op; // @[ALU.scala 35:42]
  reg [15:0] input_; // @[ALU.scala 36:42]
  reg  sourceLeftInput; // @[ALU.scala 38:32]
  reg  sourceRightInput; // @[ALU.scala 40:32]
  reg  destInput; // @[ALU.scala 41:46]
  reg [15:0] reg_0; // @[ALU.scala 43:20]
  wire [15:0] sourceLeft = ~sourceLeftInput ? $signed(input_) : $signed(reg_0); // @[ALU.scala 45:8]
  wire [15:0] sourceRight = ~sourceRightInput ? $signed(input_) : $signed(reg_0); // @[ALU.scala 47:8]
  wire  _dest_T_2 = ~destInput | op == 4'h0; // @[ALU.scala 51:25]
  wire  _result_T_54 = $signed(sourceLeft) < $signed(sourceRight); // @[ALU.scala 128:29]
  wire [15:0] _result_T_55 = $signed(sourceLeft) < $signed(sourceRight) ? $signed(sourceRight) : $signed(sourceLeft); // @[ALU.scala 128:29]
  wire [15:0] _result_T_53 = _result_T_54 ? $signed(sourceLeft) : $signed(sourceRight); // @[ALU.scala 125:29]
  wire [15:0] _GEN_17 = $signed(sourceLeft) >= $signed(sourceRight) ? $signed(16'sh100) : $signed(16'sh0); // @[ALU.scala 119:12 120:37 121:14]
  wire [15:0] _GEN_15 = $signed(sourceLeft) > $signed(sourceRight) ? $signed(16'sh100) : $signed(16'sh0); // @[ALU.scala 113:12 114:36 115:14]
  wire [15:0] _result_T_42 = 16'sh0 - $signed(sourceLeft); // @[ALU.scala 108:26]
  wire [15:0] _result_T_43 = $signed(sourceLeft) < 16'sh0 ? $signed(_result_T_42) : $signed(sourceLeft); // @[ALU.scala 108:26]
  wire [31:0] _result_mac_T_8 = $signed(sourceLeft) * $signed(sourceRight); // @[package.scala 117:18]
  wire [32:0] result_mac_4 = {{1{_result_mac_T_8[31]}},_result_mac_T_8}; // @[package.scala 117:23]
  wire [24:0] _result_adjusted_T_12 = result_mac_4[32:8]; // @[package.scala 130:26]
  wire [32:0] _result_adjustment_T_45 = $signed(result_mac_4) & 33'sh80; // @[package.scala 125:16]
  wire [8:0] result_mask1_4 = 9'sh80 - 9'sh1; // @[package.scala 120:44]
  wire [32:0] _GEN_21 = {{24{result_mask1_4[8]}},result_mask1_4}; // @[package.scala 125:44]
  wire [32:0] _result_adjustment_T_48 = $signed(result_mac_4) & $signed(_GEN_21); // @[package.scala 125:44]
  wire [32:0] _result_adjustment_T_51 = $signed(result_mac_4) & 33'sh100; // @[package.scala 125:71]
  wire  _result_adjustment_T_54 = $signed(_result_adjustment_T_45) != 33'sh0 & ($signed(_result_adjustment_T_48) != 33'sh0
     | $signed(_result_adjustment_T_51) != 33'sh0); // @[package.scala 125:34]
  wire [1:0] result_adjustment_4 = _result_adjustment_T_54 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [24:0] _GEN_22 = {{23{result_adjustment_4[1]}},result_adjustment_4}; // @[package.scala 130:42]
  wire [24:0] result_adjusted_4 = $signed(_result_adjusted_T_12) + $signed(_GEN_22); // @[package.scala 130:42]
  wire [24:0] _result_saturated_T_14 = $signed(result_adjusted_4) < -25'sh8000 ? $signed(-25'sh8000) : $signed(
    result_adjusted_4); // @[package.scala 98:26]
  wire [24:0] result_saturated_4 = $signed(result_adjusted_4) > 25'sh7fff ? $signed(25'sh7fff) : $signed(
    _result_saturated_T_14); // @[package.scala 98:8]
  wire [25:0] _result_mac_T_6 = $signed(sourceLeft) * 10'sh100; // @[package.scala 117:18]
  wire [16:0] _result_T_33 = 16'sh0 - $signed(sourceRight); // @[package.scala 171:45]
  wire [24:0] _result_mac_T_7 = {$signed(_result_T_33), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_23 = {{1{_result_mac_T_7[24]}},_result_mac_T_7}; // @[package.scala 117:23]
  wire [26:0] result_mac_3 = $signed(_result_mac_T_6) + $signed(_GEN_23); // @[package.scala 117:23]
  wire [18:0] _result_adjusted_T_9 = result_mac_3[26:8]; // @[package.scala 130:26]
  wire [26:0] _result_adjustment_T_34 = $signed(result_mac_3) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _GEN_24 = {{18{result_mask1_4[8]}},result_mask1_4}; // @[package.scala 125:44]
  wire [26:0] _result_adjustment_T_37 = $signed(result_mac_3) & $signed(_GEN_24); // @[package.scala 125:44]
  wire [26:0] _result_adjustment_T_40 = $signed(result_mac_3) & 27'sh100; // @[package.scala 125:71]
  wire  _result_adjustment_T_43 = $signed(_result_adjustment_T_34) != 27'sh0 & ($signed(_result_adjustment_T_37) != 27'sh0
     | $signed(_result_adjustment_T_40) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] result_adjustment_3 = _result_adjustment_T_43 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _GEN_25 = {{17{result_adjustment_3[1]}},result_adjustment_3}; // @[package.scala 130:42]
  wire [18:0] result_adjusted_3 = $signed(_result_adjusted_T_9) + $signed(_GEN_25); // @[package.scala 130:42]
  wire [18:0] _result_saturated_T_11 = $signed(result_adjusted_3) < -19'sh8000 ? $signed(-19'sh8000) : $signed(
    result_adjusted_3); // @[package.scala 98:26]
  wire [18:0] result_saturated_3 = $signed(result_adjusted_3) > 19'sh7fff ? $signed(19'sh7fff) : $signed(
    _result_saturated_T_11); // @[package.scala 98:8]
  wire [23:0] _result_mac_T_5 = {$signed(sourceRight), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_26 = {{2{_result_mac_T_5[23]}},_result_mac_T_5}; // @[package.scala 117:23]
  wire [26:0] result_mac_2 = $signed(_result_mac_T_6) + $signed(_GEN_26); // @[package.scala 117:23]
  wire [18:0] _result_adjusted_T_6 = result_mac_2[26:8]; // @[package.scala 130:26]
  wire [26:0] _result_adjustment_T_23 = $signed(result_mac_2) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _result_adjustment_T_26 = $signed(result_mac_2) & $signed(_GEN_24); // @[package.scala 125:44]
  wire [26:0] _result_adjustment_T_29 = $signed(result_mac_2) & 27'sh100; // @[package.scala 125:71]
  wire  _result_adjustment_T_32 = $signed(_result_adjustment_T_23) != 27'sh0 & ($signed(_result_adjustment_T_26) != 27'sh0
     | $signed(_result_adjustment_T_29) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] result_adjustment_2 = _result_adjustment_T_32 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _GEN_28 = {{17{result_adjustment_2[1]}},result_adjustment_2}; // @[package.scala 130:42]
  wire [18:0] result_adjusted_2 = $signed(_result_adjusted_T_6) + $signed(_GEN_28); // @[package.scala 130:42]
  wire [18:0] _result_saturated_T_8 = $signed(result_adjusted_2) < -19'sh8000 ? $signed(-19'sh8000) : $signed(
    result_adjusted_2); // @[package.scala 98:26]
  wire [18:0] result_saturated_2 = $signed(result_adjusted_2) > 19'sh7fff ? $signed(19'sh7fff) : $signed(
    _result_saturated_T_8); // @[package.scala 98:8]
  wire [16:0] _result_T_24 = 16'sh0 - 16'sh100; // @[package.scala 171:45]
  wire [24:0] _result_mac_T_3 = {$signed(_result_T_24), 8'h0}; // @[package.scala 117:29]
  wire [25:0] _GEN_29 = {{1{_result_mac_T_3[24]}},_result_mac_T_3}; // @[package.scala 117:23]
  wire [26:0] result_mac_1 = $signed(_result_mac_T_6) + $signed(_GEN_29); // @[package.scala 117:23]
  wire [18:0] _result_adjusted_T_3 = result_mac_1[26:8]; // @[package.scala 130:26]
  wire [26:0] _result_adjustment_T_12 = $signed(result_mac_1) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _result_adjustment_T_15 = $signed(result_mac_1) & $signed(_GEN_24); // @[package.scala 125:44]
  wire [26:0] _result_adjustment_T_18 = $signed(result_mac_1) & 27'sh100; // @[package.scala 125:71]
  wire  _result_adjustment_T_21 = $signed(_result_adjustment_T_12) != 27'sh0 & ($signed(_result_adjustment_T_15) != 27'sh0
     | $signed(_result_adjustment_T_18) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] result_adjustment_1 = _result_adjustment_T_21 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _GEN_31 = {{17{result_adjustment_1[1]}},result_adjustment_1}; // @[package.scala 130:42]
  wire [18:0] result_adjusted_1 = $signed(_result_adjusted_T_3) + $signed(_GEN_31); // @[package.scala 130:42]
  wire [18:0] _result_saturated_T_5 = $signed(result_adjusted_1) < -19'sh8000 ? $signed(-19'sh8000) : $signed(
    result_adjusted_1); // @[package.scala 98:26]
  wire [18:0] result_saturated_1 = $signed(result_adjusted_1) > 19'sh7fff ? $signed(19'sh7fff) : $signed(
    _result_saturated_T_5); // @[package.scala 98:8]
  wire [26:0] result_mac = $signed(_result_mac_T_6) + 26'sh10000; // @[package.scala 117:23]
  wire [18:0] _result_adjusted_T = result_mac[26:8]; // @[package.scala 130:26]
  wire [26:0] _result_adjustment_T_1 = $signed(result_mac) & 27'sh80; // @[package.scala 125:16]
  wire [26:0] _result_adjustment_T_4 = $signed(result_mac) & $signed(_GEN_24); // @[package.scala 125:44]
  wire [26:0] _result_adjustment_T_7 = $signed(result_mac) & 27'sh100; // @[package.scala 125:71]
  wire  _result_adjustment_T_10 = $signed(_result_adjustment_T_1) != 27'sh0 & ($signed(_result_adjustment_T_4) != 27'sh0
     | $signed(_result_adjustment_T_7) != 27'sh0); // @[package.scala 125:34]
  wire [1:0] result_adjustment = _result_adjustment_T_10 ? $signed(2'sh1) : $signed(2'sh0); // @[package.scala 124:10]
  wire [18:0] _GEN_33 = {{17{result_adjustment[1]}},result_adjustment}; // @[package.scala 130:42]
  wire [18:0] result_adjusted = $signed(_result_adjusted_T) + $signed(_GEN_33); // @[package.scala 130:42]
  wire [18:0] _result_saturated_T_2 = $signed(result_adjusted) < -19'sh8000 ? $signed(-19'sh8000) : $signed(
    result_adjusted); // @[package.scala 98:26]
  wire [18:0] result_saturated = $signed(result_adjusted) > 19'sh7fff ? $signed(19'sh7fff) : $signed(
    _result_saturated_T_2); // @[package.scala 98:8]
  wire  _T_28 = $signed(sourceLeft) >= 16'sh0 & 16'sh0 >= $signed(sourceLeft); // @[ALU.scala 132:54]
  wire  _T_29 = ~_T_28; // @[ALU.scala 131:40]
  wire  _T_34 = $signed(sourceRight) >= 16'sh0 & 16'sh0 >= $signed(sourceRight); // @[ALU.scala 132:54]
  wire  _T_35 = ~_T_34; // @[ALU.scala 131:40]
  wire [15:0] _GEN_7 = _T_29 | _T_35 ? $signed(16'sh100) : $signed(16'sh0); // @[ALU.scala 85:12 86:53 87:14]
  wire [15:0] _GEN_5 = _T_29 & _T_35 ? $signed(16'sh100) : $signed(16'sh0); // @[ALU.scala 79:12 80:53 81:14]
  wire [15:0] _GEN_3 = _T_29 ? $signed(16'sh0) : $signed(16'sh100); // @[ALU.scala 73:12 74:30 75:14]
  wire [15:0] _GEN_1 = op == 4'h1 ? $signed(16'sh0) : $signed(input_); // @[ALU.scala 62:10 64:26 65:12]
  wire [15:0] _GEN_2 = op == 4'h2 ? $signed(sourceLeft) : $signed(_GEN_1); // @[ALU.scala 67:26 68:12]
  wire [15:0] _GEN_4 = op == 4'h3 ? $signed(_GEN_3) : $signed(_GEN_2); // @[ALU.scala 72:25]
  wire [15:0] _GEN_6 = op == 4'h4 ? $signed(_GEN_5) : $signed(_GEN_4); // @[ALU.scala 78:25]
  wire [15:0] _GEN_8 = op == 4'h5 ? $signed(_GEN_7) : $signed(_GEN_6); // @[ALU.scala 84:24]
  wire [18:0] _GEN_9 = op == 4'h6 ? $signed(result_saturated) : $signed({{3{_GEN_8[15]}},_GEN_8}); // @[ALU.scala 92:31 93:12]
  wire [18:0] _GEN_10 = op == 4'h7 ? $signed(result_saturated_1) : $signed(_GEN_9); // @[ALU.scala 95:31 96:12]
  wire [18:0] _GEN_11 = op == 4'h8 ? $signed(result_saturated_2) : $signed(_GEN_10); // @[ALU.scala 98:25 99:12]
  wire [18:0] _GEN_12 = op == 4'h9 ? $signed(result_saturated_3) : $signed(_GEN_11); // @[ALU.scala 101:30 102:12]
  wire [24:0] _GEN_13 = op == 4'ha ? $signed(result_saturated_4) : $signed({{6{_GEN_12[18]}},_GEN_12}); // @[ALU.scala 104:30 105:12]
  wire [24:0] _GEN_14 = op == 4'hb ? $signed({{9{_result_T_43[15]}},_result_T_43}) : $signed(_GEN_13); // @[ALU.scala 107:25 108:12]
  wire [24:0] _GEN_16 = op == 4'hc ? $signed({{9{_GEN_15[15]}},_GEN_15}) : $signed(_GEN_14); // @[ALU.scala 112:33]
  wire [24:0] _GEN_18 = op == 4'hd ? $signed({{9{_GEN_17[15]}},_GEN_17}) : $signed(_GEN_16); // @[ALU.scala 118:38]
  wire [24:0] _GEN_19 = op == 4'he ? $signed({{9{_result_T_53[15]}},_result_T_53}) : $signed(_GEN_18); // @[ALU.scala 124:25 125:12]
  wire [24:0] _GEN_20 = op == 4'hf ? $signed({{9{_result_T_55[15]}},_result_T_55}) : $signed(_GEN_19); // @[ALU.scala 127:25 128:12]
  wire [15:0] result = _GEN_20[15:0]; // @[ALU.scala 56:20]
  reg [15:0] output_; // @[ALU.scala 57:43]
  assign io_output = output_; // @[ALU.scala 58:13]
  always @(posedge clock) begin
    op <= io_op; // @[ALU.scala 35:42]
    input_ <= io_input; // @[ALU.scala 36:42]
    sourceLeftInput <= io_sourceLeft; // @[ALU.scala 38:32]
    sourceRightInput <= io_sourceRight; // @[ALU.scala 40:32]
    destInput <= io_dest; // @[ALU.scala 41:46]
    if (reset) begin // @[ALU.scala 43:20]
      reg_0 <= 16'sh0; // @[ALU.scala 43:20]
    end else if (!(_dest_T_2)) begin // @[Demux.scala 12:16]
      reg_0 <= result; // @[Demux.scala 15:11]
    end
    output_ <= _GEN_20[15:0]; // @[ALU.scala 56:20]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  op = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  input_ = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  sourceLeftInput = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  sourceRightInput = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  destInput = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  reg_0 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  output_ = _RAND_6[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALUArray(
  input         clock,
  input         reset,
  output        io_input_ready,
  input         io_input_valid,
  input  [15:0] io_input_bits_0,
  input  [15:0] io_input_bits_1,
  input  [15:0] io_input_bits_2,
  input  [15:0] io_input_bits_3,
  input  [15:0] io_input_bits_4,
  input  [15:0] io_input_bits_5,
  input  [15:0] io_input_bits_6,
  input  [15:0] io_input_bits_7,
  input  [15:0] io_input_bits_8,
  input  [15:0] io_input_bits_9,
  input  [15:0] io_input_bits_10,
  input  [15:0] io_input_bits_11,
  input  [15:0] io_input_bits_12,
  input  [15:0] io_input_bits_13,
  input  [15:0] io_input_bits_14,
  input  [15:0] io_input_bits_15,
  input  [15:0] io_input_bits_16,
  input  [15:0] io_input_bits_17,
  input  [15:0] io_input_bits_18,
  input  [15:0] io_input_bits_19,
  input  [15:0] io_input_bits_20,
  input  [15:0] io_input_bits_21,
  input  [15:0] io_input_bits_22,
  input  [15:0] io_input_bits_23,
  input  [15:0] io_input_bits_24,
  input  [15:0] io_input_bits_25,
  input  [15:0] io_input_bits_26,
  input  [15:0] io_input_bits_27,
  input  [15:0] io_input_bits_28,
  input  [15:0] io_input_bits_29,
  input  [15:0] io_input_bits_30,
  input  [15:0] io_input_bits_31,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_0,
  output [15:0] io_output_bits_1,
  output [15:0] io_output_bits_2,
  output [15:0] io_output_bits_3,
  output [15:0] io_output_bits_4,
  output [15:0] io_output_bits_5,
  output [15:0] io_output_bits_6,
  output [15:0] io_output_bits_7,
  output [15:0] io_output_bits_8,
  output [15:0] io_output_bits_9,
  output [15:0] io_output_bits_10,
  output [15:0] io_output_bits_11,
  output [15:0] io_output_bits_12,
  output [15:0] io_output_bits_13,
  output [15:0] io_output_bits_14,
  output [15:0] io_output_bits_15,
  output [15:0] io_output_bits_16,
  output [15:0] io_output_bits_17,
  output [15:0] io_output_bits_18,
  output [15:0] io_output_bits_19,
  output [15:0] io_output_bits_20,
  output [15:0] io_output_bits_21,
  output [15:0] io_output_bits_22,
  output [15:0] io_output_bits_23,
  output [15:0] io_output_bits_24,
  output [15:0] io_output_bits_25,
  output [15:0] io_output_bits_26,
  output [15:0] io_output_bits_27,
  output [15:0] io_output_bits_28,
  output [15:0] io_output_bits_29,
  output [15:0] io_output_bits_30,
  output [15:0] io_output_bits_31,
  output        io_instruction_ready,
  input         io_instruction_valid,
  input  [3:0]  io_instruction_bits_op,
  input         io_instruction_bits_sourceLeft,
  input         io_instruction_bits_sourceRight,
  input         io_instruction_bits_dest
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  output__clock; // @[ALUArray.scala 34:22]
  wire  output__reset; // @[ALUArray.scala 34:22]
  wire  output__io_enq_ready; // @[ALUArray.scala 34:22]
  wire  output__io_enq_valid; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_0; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_1; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_2; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_3; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_4; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_5; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_6; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_7; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_8; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_9; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_10; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_11; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_12; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_13; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_14; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_15; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_16; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_17; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_18; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_19; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_20; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_21; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_22; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_23; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_24; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_25; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_26; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_27; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_28; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_29; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_30; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_enq_bits_31; // @[ALUArray.scala 34:22]
  wire  output__io_deq_ready; // @[ALUArray.scala 34:22]
  wire  output__io_deq_valid; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_0; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_1; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_2; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_3; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_4; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_5; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_6; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_7; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_8; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_9; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_10; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_11; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_12; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_13; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_14; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_15; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_16; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_17; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_18; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_19; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_20; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_21; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_22; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_23; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_24; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_25; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_26; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_27; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_28; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_29; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_30; // @[ALUArray.scala 34:22]
  wire [15:0] output__io_deq_bits_31; // @[ALUArray.scala 34:22]
  wire  m_clock; // @[ALUArray.scala 53:19]
  wire  m_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_io_input; // @[ALUArray.scala 53:19]
  wire  m_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_io_output; // @[ALUArray.scala 53:19]
  wire  m_1_clock; // @[ALUArray.scala 53:19]
  wire  m_1_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_1_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_1_io_input; // @[ALUArray.scala 53:19]
  wire  m_1_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_1_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_1_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_1_io_output; // @[ALUArray.scala 53:19]
  wire  m_2_clock; // @[ALUArray.scala 53:19]
  wire  m_2_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_2_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_2_io_input; // @[ALUArray.scala 53:19]
  wire  m_2_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_2_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_2_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_2_io_output; // @[ALUArray.scala 53:19]
  wire  m_3_clock; // @[ALUArray.scala 53:19]
  wire  m_3_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_3_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_3_io_input; // @[ALUArray.scala 53:19]
  wire  m_3_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_3_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_3_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_3_io_output; // @[ALUArray.scala 53:19]
  wire  m_4_clock; // @[ALUArray.scala 53:19]
  wire  m_4_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_4_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_4_io_input; // @[ALUArray.scala 53:19]
  wire  m_4_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_4_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_4_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_4_io_output; // @[ALUArray.scala 53:19]
  wire  m_5_clock; // @[ALUArray.scala 53:19]
  wire  m_5_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_5_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_5_io_input; // @[ALUArray.scala 53:19]
  wire  m_5_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_5_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_5_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_5_io_output; // @[ALUArray.scala 53:19]
  wire  m_6_clock; // @[ALUArray.scala 53:19]
  wire  m_6_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_6_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_6_io_input; // @[ALUArray.scala 53:19]
  wire  m_6_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_6_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_6_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_6_io_output; // @[ALUArray.scala 53:19]
  wire  m_7_clock; // @[ALUArray.scala 53:19]
  wire  m_7_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_7_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_7_io_input; // @[ALUArray.scala 53:19]
  wire  m_7_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_7_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_7_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_7_io_output; // @[ALUArray.scala 53:19]
  wire  m_8_clock; // @[ALUArray.scala 53:19]
  wire  m_8_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_8_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_8_io_input; // @[ALUArray.scala 53:19]
  wire  m_8_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_8_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_8_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_8_io_output; // @[ALUArray.scala 53:19]
  wire  m_9_clock; // @[ALUArray.scala 53:19]
  wire  m_9_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_9_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_9_io_input; // @[ALUArray.scala 53:19]
  wire  m_9_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_9_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_9_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_9_io_output; // @[ALUArray.scala 53:19]
  wire  m_10_clock; // @[ALUArray.scala 53:19]
  wire  m_10_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_10_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_10_io_input; // @[ALUArray.scala 53:19]
  wire  m_10_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_10_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_10_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_10_io_output; // @[ALUArray.scala 53:19]
  wire  m_11_clock; // @[ALUArray.scala 53:19]
  wire  m_11_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_11_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_11_io_input; // @[ALUArray.scala 53:19]
  wire  m_11_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_11_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_11_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_11_io_output; // @[ALUArray.scala 53:19]
  wire  m_12_clock; // @[ALUArray.scala 53:19]
  wire  m_12_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_12_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_12_io_input; // @[ALUArray.scala 53:19]
  wire  m_12_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_12_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_12_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_12_io_output; // @[ALUArray.scala 53:19]
  wire  m_13_clock; // @[ALUArray.scala 53:19]
  wire  m_13_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_13_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_13_io_input; // @[ALUArray.scala 53:19]
  wire  m_13_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_13_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_13_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_13_io_output; // @[ALUArray.scala 53:19]
  wire  m_14_clock; // @[ALUArray.scala 53:19]
  wire  m_14_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_14_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_14_io_input; // @[ALUArray.scala 53:19]
  wire  m_14_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_14_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_14_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_14_io_output; // @[ALUArray.scala 53:19]
  wire  m_15_clock; // @[ALUArray.scala 53:19]
  wire  m_15_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_15_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_15_io_input; // @[ALUArray.scala 53:19]
  wire  m_15_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_15_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_15_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_15_io_output; // @[ALUArray.scala 53:19]
  wire  m_16_clock; // @[ALUArray.scala 53:19]
  wire  m_16_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_16_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_16_io_input; // @[ALUArray.scala 53:19]
  wire  m_16_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_16_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_16_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_16_io_output; // @[ALUArray.scala 53:19]
  wire  m_17_clock; // @[ALUArray.scala 53:19]
  wire  m_17_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_17_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_17_io_input; // @[ALUArray.scala 53:19]
  wire  m_17_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_17_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_17_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_17_io_output; // @[ALUArray.scala 53:19]
  wire  m_18_clock; // @[ALUArray.scala 53:19]
  wire  m_18_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_18_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_18_io_input; // @[ALUArray.scala 53:19]
  wire  m_18_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_18_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_18_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_18_io_output; // @[ALUArray.scala 53:19]
  wire  m_19_clock; // @[ALUArray.scala 53:19]
  wire  m_19_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_19_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_19_io_input; // @[ALUArray.scala 53:19]
  wire  m_19_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_19_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_19_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_19_io_output; // @[ALUArray.scala 53:19]
  wire  m_20_clock; // @[ALUArray.scala 53:19]
  wire  m_20_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_20_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_20_io_input; // @[ALUArray.scala 53:19]
  wire  m_20_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_20_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_20_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_20_io_output; // @[ALUArray.scala 53:19]
  wire  m_21_clock; // @[ALUArray.scala 53:19]
  wire  m_21_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_21_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_21_io_input; // @[ALUArray.scala 53:19]
  wire  m_21_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_21_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_21_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_21_io_output; // @[ALUArray.scala 53:19]
  wire  m_22_clock; // @[ALUArray.scala 53:19]
  wire  m_22_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_22_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_22_io_input; // @[ALUArray.scala 53:19]
  wire  m_22_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_22_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_22_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_22_io_output; // @[ALUArray.scala 53:19]
  wire  m_23_clock; // @[ALUArray.scala 53:19]
  wire  m_23_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_23_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_23_io_input; // @[ALUArray.scala 53:19]
  wire  m_23_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_23_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_23_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_23_io_output; // @[ALUArray.scala 53:19]
  wire  m_24_clock; // @[ALUArray.scala 53:19]
  wire  m_24_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_24_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_24_io_input; // @[ALUArray.scala 53:19]
  wire  m_24_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_24_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_24_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_24_io_output; // @[ALUArray.scala 53:19]
  wire  m_25_clock; // @[ALUArray.scala 53:19]
  wire  m_25_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_25_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_25_io_input; // @[ALUArray.scala 53:19]
  wire  m_25_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_25_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_25_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_25_io_output; // @[ALUArray.scala 53:19]
  wire  m_26_clock; // @[ALUArray.scala 53:19]
  wire  m_26_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_26_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_26_io_input; // @[ALUArray.scala 53:19]
  wire  m_26_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_26_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_26_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_26_io_output; // @[ALUArray.scala 53:19]
  wire  m_27_clock; // @[ALUArray.scala 53:19]
  wire  m_27_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_27_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_27_io_input; // @[ALUArray.scala 53:19]
  wire  m_27_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_27_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_27_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_27_io_output; // @[ALUArray.scala 53:19]
  wire  m_28_clock; // @[ALUArray.scala 53:19]
  wire  m_28_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_28_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_28_io_input; // @[ALUArray.scala 53:19]
  wire  m_28_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_28_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_28_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_28_io_output; // @[ALUArray.scala 53:19]
  wire  m_29_clock; // @[ALUArray.scala 53:19]
  wire  m_29_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_29_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_29_io_input; // @[ALUArray.scala 53:19]
  wire  m_29_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_29_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_29_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_29_io_output; // @[ALUArray.scala 53:19]
  wire  m_30_clock; // @[ALUArray.scala 53:19]
  wire  m_30_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_30_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_30_io_input; // @[ALUArray.scala 53:19]
  wire  m_30_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_30_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_30_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_30_io_output; // @[ALUArray.scala 53:19]
  wire  m_31_clock; // @[ALUArray.scala 53:19]
  wire  m_31_reset; // @[ALUArray.scala 53:19]
  wire [3:0] m_31_io_op; // @[ALUArray.scala 53:19]
  wire [15:0] m_31_io_input; // @[ALUArray.scala 53:19]
  wire  m_31_io_sourceLeft; // @[ALUArray.scala 53:19]
  wire  m_31_io_sourceRight; // @[ALUArray.scala 53:19]
  wire  m_31_io_dest; // @[ALUArray.scala 53:19]
  wire [15:0] m_31_io_output; // @[ALUArray.scala 53:19]
  wire  _inputNotNeeded_T_11 = io_instruction_bits_op == 4'h2 & io_instruction_bits_op == 4'h3 & io_instruction_bits_op
     == 4'h6 & io_instruction_bits_op == 4'h7 & io_instruction_bits_op == 4'hb; // @[Op.scala 40:39]
  wire  _inputNotNeeded_T_13 = _inputNotNeeded_T_11 & io_instruction_bits_sourceLeft; // @[ALUArray.scala 41:9]
  wire  _inputNotNeeded_T_14 = io_instruction_bits_op == 4'h0 | io_instruction_bits_op == 4'h1 | _inputNotNeeded_T_13; // @[ALUArray.scala 38:76]
  wire  _inputNotNeeded_T_17 = io_instruction_bits_sourceLeft & io_instruction_bits_sourceRight; // @[ALUArray.scala 42:44]
  wire  inputNotNeeded = _inputNotNeeded_T_14 | _inputNotNeeded_T_17; // @[ALUArray.scala 41:49]
  wire  inputNeeded = ~inputNotNeeded; // @[ALUArray.scala 43:21]
  wire  _io_instruction_ready_T_1 = io_input_valid | ~inputNeeded; // @[ALUArray.scala 46:38]
  wire  _output_io_enq_valid_T_2 = _io_instruction_ready_T_1 & io_instruction_valid; // @[ALUArray.scala 48:35]
  reg  output_io_enq_valid_sr_0; // @[ShiftRegister.scala 10:22]
  reg  output_io_enq_valid_sr_1; // @[ShiftRegister.scala 10:22]
  wire  _m_io_op_T = io_instruction_ready & io_instruction_valid; // @[ALUArray.scala 63:25]
  Queue_17 output_ ( // @[ALUArray.scala 34:22]
    .clock(output__clock),
    .reset(output__reset),
    .io_enq_ready(output__io_enq_ready),
    .io_enq_valid(output__io_enq_valid),
    .io_enq_bits_0(output__io_enq_bits_0),
    .io_enq_bits_1(output__io_enq_bits_1),
    .io_enq_bits_2(output__io_enq_bits_2),
    .io_enq_bits_3(output__io_enq_bits_3),
    .io_enq_bits_4(output__io_enq_bits_4),
    .io_enq_bits_5(output__io_enq_bits_5),
    .io_enq_bits_6(output__io_enq_bits_6),
    .io_enq_bits_7(output__io_enq_bits_7),
    .io_enq_bits_8(output__io_enq_bits_8),
    .io_enq_bits_9(output__io_enq_bits_9),
    .io_enq_bits_10(output__io_enq_bits_10),
    .io_enq_bits_11(output__io_enq_bits_11),
    .io_enq_bits_12(output__io_enq_bits_12),
    .io_enq_bits_13(output__io_enq_bits_13),
    .io_enq_bits_14(output__io_enq_bits_14),
    .io_enq_bits_15(output__io_enq_bits_15),
    .io_enq_bits_16(output__io_enq_bits_16),
    .io_enq_bits_17(output__io_enq_bits_17),
    .io_enq_bits_18(output__io_enq_bits_18),
    .io_enq_bits_19(output__io_enq_bits_19),
    .io_enq_bits_20(output__io_enq_bits_20),
    .io_enq_bits_21(output__io_enq_bits_21),
    .io_enq_bits_22(output__io_enq_bits_22),
    .io_enq_bits_23(output__io_enq_bits_23),
    .io_enq_bits_24(output__io_enq_bits_24),
    .io_enq_bits_25(output__io_enq_bits_25),
    .io_enq_bits_26(output__io_enq_bits_26),
    .io_enq_bits_27(output__io_enq_bits_27),
    .io_enq_bits_28(output__io_enq_bits_28),
    .io_enq_bits_29(output__io_enq_bits_29),
    .io_enq_bits_30(output__io_enq_bits_30),
    .io_enq_bits_31(output__io_enq_bits_31),
    .io_deq_ready(output__io_deq_ready),
    .io_deq_valid(output__io_deq_valid),
    .io_deq_bits_0(output__io_deq_bits_0),
    .io_deq_bits_1(output__io_deq_bits_1),
    .io_deq_bits_2(output__io_deq_bits_2),
    .io_deq_bits_3(output__io_deq_bits_3),
    .io_deq_bits_4(output__io_deq_bits_4),
    .io_deq_bits_5(output__io_deq_bits_5),
    .io_deq_bits_6(output__io_deq_bits_6),
    .io_deq_bits_7(output__io_deq_bits_7),
    .io_deq_bits_8(output__io_deq_bits_8),
    .io_deq_bits_9(output__io_deq_bits_9),
    .io_deq_bits_10(output__io_deq_bits_10),
    .io_deq_bits_11(output__io_deq_bits_11),
    .io_deq_bits_12(output__io_deq_bits_12),
    .io_deq_bits_13(output__io_deq_bits_13),
    .io_deq_bits_14(output__io_deq_bits_14),
    .io_deq_bits_15(output__io_deq_bits_15),
    .io_deq_bits_16(output__io_deq_bits_16),
    .io_deq_bits_17(output__io_deq_bits_17),
    .io_deq_bits_18(output__io_deq_bits_18),
    .io_deq_bits_19(output__io_deq_bits_19),
    .io_deq_bits_20(output__io_deq_bits_20),
    .io_deq_bits_21(output__io_deq_bits_21),
    .io_deq_bits_22(output__io_deq_bits_22),
    .io_deq_bits_23(output__io_deq_bits_23),
    .io_deq_bits_24(output__io_deq_bits_24),
    .io_deq_bits_25(output__io_deq_bits_25),
    .io_deq_bits_26(output__io_deq_bits_26),
    .io_deq_bits_27(output__io_deq_bits_27),
    .io_deq_bits_28(output__io_deq_bits_28),
    .io_deq_bits_29(output__io_deq_bits_29),
    .io_deq_bits_30(output__io_deq_bits_30),
    .io_deq_bits_31(output__io_deq_bits_31)
  );
  ALU m ( // @[ALUArray.scala 53:19]
    .clock(m_clock),
    .reset(m_reset),
    .io_op(m_io_op),
    .io_input(m_io_input),
    .io_sourceLeft(m_io_sourceLeft),
    .io_sourceRight(m_io_sourceRight),
    .io_dest(m_io_dest),
    .io_output(m_io_output)
  );
  ALU m_1 ( // @[ALUArray.scala 53:19]
    .clock(m_1_clock),
    .reset(m_1_reset),
    .io_op(m_1_io_op),
    .io_input(m_1_io_input),
    .io_sourceLeft(m_1_io_sourceLeft),
    .io_sourceRight(m_1_io_sourceRight),
    .io_dest(m_1_io_dest),
    .io_output(m_1_io_output)
  );
  ALU m_2 ( // @[ALUArray.scala 53:19]
    .clock(m_2_clock),
    .reset(m_2_reset),
    .io_op(m_2_io_op),
    .io_input(m_2_io_input),
    .io_sourceLeft(m_2_io_sourceLeft),
    .io_sourceRight(m_2_io_sourceRight),
    .io_dest(m_2_io_dest),
    .io_output(m_2_io_output)
  );
  ALU m_3 ( // @[ALUArray.scala 53:19]
    .clock(m_3_clock),
    .reset(m_3_reset),
    .io_op(m_3_io_op),
    .io_input(m_3_io_input),
    .io_sourceLeft(m_3_io_sourceLeft),
    .io_sourceRight(m_3_io_sourceRight),
    .io_dest(m_3_io_dest),
    .io_output(m_3_io_output)
  );
  ALU m_4 ( // @[ALUArray.scala 53:19]
    .clock(m_4_clock),
    .reset(m_4_reset),
    .io_op(m_4_io_op),
    .io_input(m_4_io_input),
    .io_sourceLeft(m_4_io_sourceLeft),
    .io_sourceRight(m_4_io_sourceRight),
    .io_dest(m_4_io_dest),
    .io_output(m_4_io_output)
  );
  ALU m_5 ( // @[ALUArray.scala 53:19]
    .clock(m_5_clock),
    .reset(m_5_reset),
    .io_op(m_5_io_op),
    .io_input(m_5_io_input),
    .io_sourceLeft(m_5_io_sourceLeft),
    .io_sourceRight(m_5_io_sourceRight),
    .io_dest(m_5_io_dest),
    .io_output(m_5_io_output)
  );
  ALU m_6 ( // @[ALUArray.scala 53:19]
    .clock(m_6_clock),
    .reset(m_6_reset),
    .io_op(m_6_io_op),
    .io_input(m_6_io_input),
    .io_sourceLeft(m_6_io_sourceLeft),
    .io_sourceRight(m_6_io_sourceRight),
    .io_dest(m_6_io_dest),
    .io_output(m_6_io_output)
  );
  ALU m_7 ( // @[ALUArray.scala 53:19]
    .clock(m_7_clock),
    .reset(m_7_reset),
    .io_op(m_7_io_op),
    .io_input(m_7_io_input),
    .io_sourceLeft(m_7_io_sourceLeft),
    .io_sourceRight(m_7_io_sourceRight),
    .io_dest(m_7_io_dest),
    .io_output(m_7_io_output)
  );
  ALU m_8 ( // @[ALUArray.scala 53:19]
    .clock(m_8_clock),
    .reset(m_8_reset),
    .io_op(m_8_io_op),
    .io_input(m_8_io_input),
    .io_sourceLeft(m_8_io_sourceLeft),
    .io_sourceRight(m_8_io_sourceRight),
    .io_dest(m_8_io_dest),
    .io_output(m_8_io_output)
  );
  ALU m_9 ( // @[ALUArray.scala 53:19]
    .clock(m_9_clock),
    .reset(m_9_reset),
    .io_op(m_9_io_op),
    .io_input(m_9_io_input),
    .io_sourceLeft(m_9_io_sourceLeft),
    .io_sourceRight(m_9_io_sourceRight),
    .io_dest(m_9_io_dest),
    .io_output(m_9_io_output)
  );
  ALU m_10 ( // @[ALUArray.scala 53:19]
    .clock(m_10_clock),
    .reset(m_10_reset),
    .io_op(m_10_io_op),
    .io_input(m_10_io_input),
    .io_sourceLeft(m_10_io_sourceLeft),
    .io_sourceRight(m_10_io_sourceRight),
    .io_dest(m_10_io_dest),
    .io_output(m_10_io_output)
  );
  ALU m_11 ( // @[ALUArray.scala 53:19]
    .clock(m_11_clock),
    .reset(m_11_reset),
    .io_op(m_11_io_op),
    .io_input(m_11_io_input),
    .io_sourceLeft(m_11_io_sourceLeft),
    .io_sourceRight(m_11_io_sourceRight),
    .io_dest(m_11_io_dest),
    .io_output(m_11_io_output)
  );
  ALU m_12 ( // @[ALUArray.scala 53:19]
    .clock(m_12_clock),
    .reset(m_12_reset),
    .io_op(m_12_io_op),
    .io_input(m_12_io_input),
    .io_sourceLeft(m_12_io_sourceLeft),
    .io_sourceRight(m_12_io_sourceRight),
    .io_dest(m_12_io_dest),
    .io_output(m_12_io_output)
  );
  ALU m_13 ( // @[ALUArray.scala 53:19]
    .clock(m_13_clock),
    .reset(m_13_reset),
    .io_op(m_13_io_op),
    .io_input(m_13_io_input),
    .io_sourceLeft(m_13_io_sourceLeft),
    .io_sourceRight(m_13_io_sourceRight),
    .io_dest(m_13_io_dest),
    .io_output(m_13_io_output)
  );
  ALU m_14 ( // @[ALUArray.scala 53:19]
    .clock(m_14_clock),
    .reset(m_14_reset),
    .io_op(m_14_io_op),
    .io_input(m_14_io_input),
    .io_sourceLeft(m_14_io_sourceLeft),
    .io_sourceRight(m_14_io_sourceRight),
    .io_dest(m_14_io_dest),
    .io_output(m_14_io_output)
  );
  ALU m_15 ( // @[ALUArray.scala 53:19]
    .clock(m_15_clock),
    .reset(m_15_reset),
    .io_op(m_15_io_op),
    .io_input(m_15_io_input),
    .io_sourceLeft(m_15_io_sourceLeft),
    .io_sourceRight(m_15_io_sourceRight),
    .io_dest(m_15_io_dest),
    .io_output(m_15_io_output)
  );
  ALU m_16 ( // @[ALUArray.scala 53:19]
    .clock(m_16_clock),
    .reset(m_16_reset),
    .io_op(m_16_io_op),
    .io_input(m_16_io_input),
    .io_sourceLeft(m_16_io_sourceLeft),
    .io_sourceRight(m_16_io_sourceRight),
    .io_dest(m_16_io_dest),
    .io_output(m_16_io_output)
  );
  ALU m_17 ( // @[ALUArray.scala 53:19]
    .clock(m_17_clock),
    .reset(m_17_reset),
    .io_op(m_17_io_op),
    .io_input(m_17_io_input),
    .io_sourceLeft(m_17_io_sourceLeft),
    .io_sourceRight(m_17_io_sourceRight),
    .io_dest(m_17_io_dest),
    .io_output(m_17_io_output)
  );
  ALU m_18 ( // @[ALUArray.scala 53:19]
    .clock(m_18_clock),
    .reset(m_18_reset),
    .io_op(m_18_io_op),
    .io_input(m_18_io_input),
    .io_sourceLeft(m_18_io_sourceLeft),
    .io_sourceRight(m_18_io_sourceRight),
    .io_dest(m_18_io_dest),
    .io_output(m_18_io_output)
  );
  ALU m_19 ( // @[ALUArray.scala 53:19]
    .clock(m_19_clock),
    .reset(m_19_reset),
    .io_op(m_19_io_op),
    .io_input(m_19_io_input),
    .io_sourceLeft(m_19_io_sourceLeft),
    .io_sourceRight(m_19_io_sourceRight),
    .io_dest(m_19_io_dest),
    .io_output(m_19_io_output)
  );
  ALU m_20 ( // @[ALUArray.scala 53:19]
    .clock(m_20_clock),
    .reset(m_20_reset),
    .io_op(m_20_io_op),
    .io_input(m_20_io_input),
    .io_sourceLeft(m_20_io_sourceLeft),
    .io_sourceRight(m_20_io_sourceRight),
    .io_dest(m_20_io_dest),
    .io_output(m_20_io_output)
  );
  ALU m_21 ( // @[ALUArray.scala 53:19]
    .clock(m_21_clock),
    .reset(m_21_reset),
    .io_op(m_21_io_op),
    .io_input(m_21_io_input),
    .io_sourceLeft(m_21_io_sourceLeft),
    .io_sourceRight(m_21_io_sourceRight),
    .io_dest(m_21_io_dest),
    .io_output(m_21_io_output)
  );
  ALU m_22 ( // @[ALUArray.scala 53:19]
    .clock(m_22_clock),
    .reset(m_22_reset),
    .io_op(m_22_io_op),
    .io_input(m_22_io_input),
    .io_sourceLeft(m_22_io_sourceLeft),
    .io_sourceRight(m_22_io_sourceRight),
    .io_dest(m_22_io_dest),
    .io_output(m_22_io_output)
  );
  ALU m_23 ( // @[ALUArray.scala 53:19]
    .clock(m_23_clock),
    .reset(m_23_reset),
    .io_op(m_23_io_op),
    .io_input(m_23_io_input),
    .io_sourceLeft(m_23_io_sourceLeft),
    .io_sourceRight(m_23_io_sourceRight),
    .io_dest(m_23_io_dest),
    .io_output(m_23_io_output)
  );
  ALU m_24 ( // @[ALUArray.scala 53:19]
    .clock(m_24_clock),
    .reset(m_24_reset),
    .io_op(m_24_io_op),
    .io_input(m_24_io_input),
    .io_sourceLeft(m_24_io_sourceLeft),
    .io_sourceRight(m_24_io_sourceRight),
    .io_dest(m_24_io_dest),
    .io_output(m_24_io_output)
  );
  ALU m_25 ( // @[ALUArray.scala 53:19]
    .clock(m_25_clock),
    .reset(m_25_reset),
    .io_op(m_25_io_op),
    .io_input(m_25_io_input),
    .io_sourceLeft(m_25_io_sourceLeft),
    .io_sourceRight(m_25_io_sourceRight),
    .io_dest(m_25_io_dest),
    .io_output(m_25_io_output)
  );
  ALU m_26 ( // @[ALUArray.scala 53:19]
    .clock(m_26_clock),
    .reset(m_26_reset),
    .io_op(m_26_io_op),
    .io_input(m_26_io_input),
    .io_sourceLeft(m_26_io_sourceLeft),
    .io_sourceRight(m_26_io_sourceRight),
    .io_dest(m_26_io_dest),
    .io_output(m_26_io_output)
  );
  ALU m_27 ( // @[ALUArray.scala 53:19]
    .clock(m_27_clock),
    .reset(m_27_reset),
    .io_op(m_27_io_op),
    .io_input(m_27_io_input),
    .io_sourceLeft(m_27_io_sourceLeft),
    .io_sourceRight(m_27_io_sourceRight),
    .io_dest(m_27_io_dest),
    .io_output(m_27_io_output)
  );
  ALU m_28 ( // @[ALUArray.scala 53:19]
    .clock(m_28_clock),
    .reset(m_28_reset),
    .io_op(m_28_io_op),
    .io_input(m_28_io_input),
    .io_sourceLeft(m_28_io_sourceLeft),
    .io_sourceRight(m_28_io_sourceRight),
    .io_dest(m_28_io_dest),
    .io_output(m_28_io_output)
  );
  ALU m_29 ( // @[ALUArray.scala 53:19]
    .clock(m_29_clock),
    .reset(m_29_reset),
    .io_op(m_29_io_op),
    .io_input(m_29_io_input),
    .io_sourceLeft(m_29_io_sourceLeft),
    .io_sourceRight(m_29_io_sourceRight),
    .io_dest(m_29_io_dest),
    .io_output(m_29_io_output)
  );
  ALU m_30 ( // @[ALUArray.scala 53:19]
    .clock(m_30_clock),
    .reset(m_30_reset),
    .io_op(m_30_io_op),
    .io_input(m_30_io_input),
    .io_sourceLeft(m_30_io_sourceLeft),
    .io_sourceRight(m_30_io_sourceRight),
    .io_dest(m_30_io_dest),
    .io_output(m_30_io_output)
  );
  ALU m_31 ( // @[ALUArray.scala 53:19]
    .clock(m_31_clock),
    .reset(m_31_reset),
    .io_op(m_31_io_op),
    .io_input(m_31_io_input),
    .io_sourceLeft(m_31_io_sourceLeft),
    .io_sourceRight(m_31_io_sourceRight),
    .io_dest(m_31_io_dest),
    .io_output(m_31_io_output)
  );
  assign io_input_ready = output__io_enq_ready & io_instruction_valid & inputNeeded; // @[ALUArray.scala 45:59]
  assign io_output_valid = output__io_deq_valid; // @[ALUArray.scala 35:13]
  assign io_output_bits_0 = output__io_deq_bits_0; // @[ALUArray.scala 35:13]
  assign io_output_bits_1 = output__io_deq_bits_1; // @[ALUArray.scala 35:13]
  assign io_output_bits_2 = output__io_deq_bits_2; // @[ALUArray.scala 35:13]
  assign io_output_bits_3 = output__io_deq_bits_3; // @[ALUArray.scala 35:13]
  assign io_output_bits_4 = output__io_deq_bits_4; // @[ALUArray.scala 35:13]
  assign io_output_bits_5 = output__io_deq_bits_5; // @[ALUArray.scala 35:13]
  assign io_output_bits_6 = output__io_deq_bits_6; // @[ALUArray.scala 35:13]
  assign io_output_bits_7 = output__io_deq_bits_7; // @[ALUArray.scala 35:13]
  assign io_output_bits_8 = output__io_deq_bits_8; // @[ALUArray.scala 35:13]
  assign io_output_bits_9 = output__io_deq_bits_9; // @[ALUArray.scala 35:13]
  assign io_output_bits_10 = output__io_deq_bits_10; // @[ALUArray.scala 35:13]
  assign io_output_bits_11 = output__io_deq_bits_11; // @[ALUArray.scala 35:13]
  assign io_output_bits_12 = output__io_deq_bits_12; // @[ALUArray.scala 35:13]
  assign io_output_bits_13 = output__io_deq_bits_13; // @[ALUArray.scala 35:13]
  assign io_output_bits_14 = output__io_deq_bits_14; // @[ALUArray.scala 35:13]
  assign io_output_bits_15 = output__io_deq_bits_15; // @[ALUArray.scala 35:13]
  assign io_output_bits_16 = output__io_deq_bits_16; // @[ALUArray.scala 35:13]
  assign io_output_bits_17 = output__io_deq_bits_17; // @[ALUArray.scala 35:13]
  assign io_output_bits_18 = output__io_deq_bits_18; // @[ALUArray.scala 35:13]
  assign io_output_bits_19 = output__io_deq_bits_19; // @[ALUArray.scala 35:13]
  assign io_output_bits_20 = output__io_deq_bits_20; // @[ALUArray.scala 35:13]
  assign io_output_bits_21 = output__io_deq_bits_21; // @[ALUArray.scala 35:13]
  assign io_output_bits_22 = output__io_deq_bits_22; // @[ALUArray.scala 35:13]
  assign io_output_bits_23 = output__io_deq_bits_23; // @[ALUArray.scala 35:13]
  assign io_output_bits_24 = output__io_deq_bits_24; // @[ALUArray.scala 35:13]
  assign io_output_bits_25 = output__io_deq_bits_25; // @[ALUArray.scala 35:13]
  assign io_output_bits_26 = output__io_deq_bits_26; // @[ALUArray.scala 35:13]
  assign io_output_bits_27 = output__io_deq_bits_27; // @[ALUArray.scala 35:13]
  assign io_output_bits_28 = output__io_deq_bits_28; // @[ALUArray.scala 35:13]
  assign io_output_bits_29 = output__io_deq_bits_29; // @[ALUArray.scala 35:13]
  assign io_output_bits_30 = output__io_deq_bits_30; // @[ALUArray.scala 35:13]
  assign io_output_bits_31 = output__io_deq_bits_31; // @[ALUArray.scala 35:13]
  assign io_instruction_ready = (io_input_valid | ~inputNeeded) & output__io_enq_ready; // @[ALUArray.scala 46:55]
  assign output__clock = clock;
  assign output__reset = reset;
  assign output__io_enq_valid = output_io_enq_valid_sr_1; // @[ALUArray.scala 47:23]
  assign output__io_enq_bits_0 = m_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_1 = m_1_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_2 = m_2_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_3 = m_3_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_4 = m_4_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_5 = m_5_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_6 = m_6_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_7 = m_7_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_8 = m_8_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_9 = m_9_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_10 = m_10_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_11 = m_11_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_12 = m_12_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_13 = m_13_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_14 = m_14_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_15 = m_15_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_16 = m_16_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_17 = m_17_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_18 = m_18_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_19 = m_19_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_20 = m_20_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_21 = m_21_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_22 = m_22_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_23 = m_23_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_24 = m_24_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_25 = m_25_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_26 = m_26_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_27 = m_27_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_28 = m_28_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_29 = m_29_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_30 = m_30_io_output; // @[ALUArray.scala 71:27]
  assign output__io_enq_bits_31 = m_31_io_output; // @[ALUArray.scala 71:27]
  assign output__io_deq_ready = io_output_ready; // @[ALUArray.scala 35:13]
  assign m_clock = clock;
  assign m_reset = reset;
  assign m_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_io_input = io_input_bits_0; // @[ALUArray.scala 70:16]
  assign m_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_1_clock = clock;
  assign m_1_reset = reset;
  assign m_1_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_1_io_input = io_input_bits_1; // @[ALUArray.scala 70:16]
  assign m_1_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_1_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_1_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_2_clock = clock;
  assign m_2_reset = reset;
  assign m_2_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_2_io_input = io_input_bits_2; // @[ALUArray.scala 70:16]
  assign m_2_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_2_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_2_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_3_clock = clock;
  assign m_3_reset = reset;
  assign m_3_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_3_io_input = io_input_bits_3; // @[ALUArray.scala 70:16]
  assign m_3_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_3_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_3_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_4_clock = clock;
  assign m_4_reset = reset;
  assign m_4_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_4_io_input = io_input_bits_4; // @[ALUArray.scala 70:16]
  assign m_4_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_4_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_4_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_5_clock = clock;
  assign m_5_reset = reset;
  assign m_5_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_5_io_input = io_input_bits_5; // @[ALUArray.scala 70:16]
  assign m_5_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_5_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_5_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_6_clock = clock;
  assign m_6_reset = reset;
  assign m_6_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_6_io_input = io_input_bits_6; // @[ALUArray.scala 70:16]
  assign m_6_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_6_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_6_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_7_clock = clock;
  assign m_7_reset = reset;
  assign m_7_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_7_io_input = io_input_bits_7; // @[ALUArray.scala 70:16]
  assign m_7_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_7_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_7_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_8_clock = clock;
  assign m_8_reset = reset;
  assign m_8_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_8_io_input = io_input_bits_8; // @[ALUArray.scala 70:16]
  assign m_8_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_8_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_8_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_9_clock = clock;
  assign m_9_reset = reset;
  assign m_9_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_9_io_input = io_input_bits_9; // @[ALUArray.scala 70:16]
  assign m_9_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_9_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_9_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_10_clock = clock;
  assign m_10_reset = reset;
  assign m_10_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_10_io_input = io_input_bits_10; // @[ALUArray.scala 70:16]
  assign m_10_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_10_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_10_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_11_clock = clock;
  assign m_11_reset = reset;
  assign m_11_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_11_io_input = io_input_bits_11; // @[ALUArray.scala 70:16]
  assign m_11_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_11_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_11_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_12_clock = clock;
  assign m_12_reset = reset;
  assign m_12_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_12_io_input = io_input_bits_12; // @[ALUArray.scala 70:16]
  assign m_12_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_12_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_12_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_13_clock = clock;
  assign m_13_reset = reset;
  assign m_13_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_13_io_input = io_input_bits_13; // @[ALUArray.scala 70:16]
  assign m_13_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_13_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_13_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_14_clock = clock;
  assign m_14_reset = reset;
  assign m_14_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_14_io_input = io_input_bits_14; // @[ALUArray.scala 70:16]
  assign m_14_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_14_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_14_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_15_clock = clock;
  assign m_15_reset = reset;
  assign m_15_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_15_io_input = io_input_bits_15; // @[ALUArray.scala 70:16]
  assign m_15_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_15_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_15_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_16_clock = clock;
  assign m_16_reset = reset;
  assign m_16_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_16_io_input = io_input_bits_16; // @[ALUArray.scala 70:16]
  assign m_16_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_16_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_16_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_17_clock = clock;
  assign m_17_reset = reset;
  assign m_17_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_17_io_input = io_input_bits_17; // @[ALUArray.scala 70:16]
  assign m_17_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_17_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_17_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_18_clock = clock;
  assign m_18_reset = reset;
  assign m_18_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_18_io_input = io_input_bits_18; // @[ALUArray.scala 70:16]
  assign m_18_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_18_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_18_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_19_clock = clock;
  assign m_19_reset = reset;
  assign m_19_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_19_io_input = io_input_bits_19; // @[ALUArray.scala 70:16]
  assign m_19_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_19_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_19_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_20_clock = clock;
  assign m_20_reset = reset;
  assign m_20_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_20_io_input = io_input_bits_20; // @[ALUArray.scala 70:16]
  assign m_20_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_20_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_20_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_21_clock = clock;
  assign m_21_reset = reset;
  assign m_21_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_21_io_input = io_input_bits_21; // @[ALUArray.scala 70:16]
  assign m_21_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_21_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_21_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_22_clock = clock;
  assign m_22_reset = reset;
  assign m_22_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_22_io_input = io_input_bits_22; // @[ALUArray.scala 70:16]
  assign m_22_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_22_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_22_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_23_clock = clock;
  assign m_23_reset = reset;
  assign m_23_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_23_io_input = io_input_bits_23; // @[ALUArray.scala 70:16]
  assign m_23_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_23_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_23_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_24_clock = clock;
  assign m_24_reset = reset;
  assign m_24_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_24_io_input = io_input_bits_24; // @[ALUArray.scala 70:16]
  assign m_24_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_24_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_24_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_25_clock = clock;
  assign m_25_reset = reset;
  assign m_25_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_25_io_input = io_input_bits_25; // @[ALUArray.scala 70:16]
  assign m_25_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_25_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_25_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_26_clock = clock;
  assign m_26_reset = reset;
  assign m_26_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_26_io_input = io_input_bits_26; // @[ALUArray.scala 70:16]
  assign m_26_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_26_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_26_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_27_clock = clock;
  assign m_27_reset = reset;
  assign m_27_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_27_io_input = io_input_bits_27; // @[ALUArray.scala 70:16]
  assign m_27_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_27_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_27_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_28_clock = clock;
  assign m_28_reset = reset;
  assign m_28_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_28_io_input = io_input_bits_28; // @[ALUArray.scala 70:16]
  assign m_28_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_28_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_28_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_29_clock = clock;
  assign m_29_reset = reset;
  assign m_29_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_29_io_input = io_input_bits_29; // @[ALUArray.scala 70:16]
  assign m_29_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_29_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_29_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_30_clock = clock;
  assign m_30_reset = reset;
  assign m_30_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_30_io_input = io_input_bits_30; // @[ALUArray.scala 70:16]
  assign m_30_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_30_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_30_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  assign m_31_clock = clock;
  assign m_31_reset = reset;
  assign m_31_io_op = _m_io_op_T ? io_instruction_bits_op : 4'h0; // @[ALUArray.scala 62:19]
  assign m_31_io_input = io_input_bits_31; // @[ALUArray.scala 70:16]
  assign m_31_io_sourceLeft = io_instruction_bits_sourceLeft; // @[ALUArray.scala 67:21]
  assign m_31_io_sourceRight = io_instruction_bits_sourceRight; // @[ALUArray.scala 68:22]
  assign m_31_io_dest = io_instruction_bits_dest; // @[ALUArray.scala 69:15]
  always @(posedge clock) begin
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_0 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_0 <= _output_io_enq_valid_T_2; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_1 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_1 <= output_io_enq_valid_sr_0; // @[ShiftRegister.scala 13:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  output_io_enq_valid_sr_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  output_io_enq_valid_sr_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AccumulatorWithALUArray(
  input         clock,
  input         reset,
  output        io_input_ready,
  input         io_input_valid,
  input  [15:0] io_input_bits_0,
  input  [15:0] io_input_bits_1,
  input  [15:0] io_input_bits_2,
  input  [15:0] io_input_bits_3,
  input  [15:0] io_input_bits_4,
  input  [15:0] io_input_bits_5,
  input  [15:0] io_input_bits_6,
  input  [15:0] io_input_bits_7,
  input  [15:0] io_input_bits_8,
  input  [15:0] io_input_bits_9,
  input  [15:0] io_input_bits_10,
  input  [15:0] io_input_bits_11,
  input  [15:0] io_input_bits_12,
  input  [15:0] io_input_bits_13,
  input  [15:0] io_input_bits_14,
  input  [15:0] io_input_bits_15,
  input  [15:0] io_input_bits_16,
  input  [15:0] io_input_bits_17,
  input  [15:0] io_input_bits_18,
  input  [15:0] io_input_bits_19,
  input  [15:0] io_input_bits_20,
  input  [15:0] io_input_bits_21,
  input  [15:0] io_input_bits_22,
  input  [15:0] io_input_bits_23,
  input  [15:0] io_input_bits_24,
  input  [15:0] io_input_bits_25,
  input  [15:0] io_input_bits_26,
  input  [15:0] io_input_bits_27,
  input  [15:0] io_input_bits_28,
  input  [15:0] io_input_bits_29,
  input  [15:0] io_input_bits_30,
  input  [15:0] io_input_bits_31,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_0,
  output [15:0] io_output_bits_1,
  output [15:0] io_output_bits_2,
  output [15:0] io_output_bits_3,
  output [15:0] io_output_bits_4,
  output [15:0] io_output_bits_5,
  output [15:0] io_output_bits_6,
  output [15:0] io_output_bits_7,
  output [15:0] io_output_bits_8,
  output [15:0] io_output_bits_9,
  output [15:0] io_output_bits_10,
  output [15:0] io_output_bits_11,
  output [15:0] io_output_bits_12,
  output [15:0] io_output_bits_13,
  output [15:0] io_output_bits_14,
  output [15:0] io_output_bits_15,
  output [15:0] io_output_bits_16,
  output [15:0] io_output_bits_17,
  output [15:0] io_output_bits_18,
  output [15:0] io_output_bits_19,
  output [15:0] io_output_bits_20,
  output [15:0] io_output_bits_21,
  output [15:0] io_output_bits_22,
  output [15:0] io_output_bits_23,
  output [15:0] io_output_bits_24,
  output [15:0] io_output_bits_25,
  output [15:0] io_output_bits_26,
  output [15:0] io_output_bits_27,
  output [15:0] io_output_bits_28,
  output [15:0] io_output_bits_29,
  output [15:0] io_output_bits_30,
  output [15:0] io_output_bits_31,
  output        io_control_ready,
  input         io_control_valid,
  input  [3:0]  io_control_bits_instruction_op,
  input         io_control_bits_instruction_sourceLeft,
  input         io_control_bits_instruction_sourceRight,
  input         io_control_bits_instruction_dest,
  input  [11:0] io_control_bits_readAddress,
  input  [11:0] io_control_bits_writeAddress,
  input         io_control_bits_accumulate,
  input         io_control_bits_write,
  input         io_control_bits_read,
  input         io_tracepoint,
  input  [31:0] io_programCounter
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  acc_clock; // @[AccumulatorWithALUArray.scala 44:19]
  wire  acc_reset; // @[AccumulatorWithALUArray.scala 44:19]
  wire  acc_io_input_ready; // @[AccumulatorWithALUArray.scala 44:19]
  wire  acc_io_input_valid; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_0; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_1; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_2; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_3; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_4; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_5; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_6; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_7; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_8; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_9; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_10; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_11; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_12; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_13; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_14; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_15; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_16; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_17; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_18; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_19; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_20; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_21; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_22; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_23; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_24; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_25; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_26; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_27; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_28; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_29; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_30; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_input_bits_31; // @[AccumulatorWithALUArray.scala 44:19]
  wire  acc_io_output_ready; // @[AccumulatorWithALUArray.scala 44:19]
  wire  acc_io_output_valid; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_0; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_1; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_2; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_3; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_4; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_5; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_6; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_7; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_8; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_9; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_10; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_11; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_12; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_13; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_14; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_15; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_16; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_17; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_18; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_19; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_20; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_21; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_22; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_23; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_24; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_25; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_26; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_27; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_28; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_29; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_30; // @[AccumulatorWithALUArray.scala 44:19]
  wire [15:0] acc_io_output_bits_31; // @[AccumulatorWithALUArray.scala 44:19]
  wire  acc_io_control_ready; // @[AccumulatorWithALUArray.scala 44:19]
  wire  acc_io_control_valid; // @[AccumulatorWithALUArray.scala 44:19]
  wire [11:0] acc_io_control_bits_address; // @[AccumulatorWithALUArray.scala 44:19]
  wire  acc_io_control_bits_accumulate; // @[AccumulatorWithALUArray.scala 44:19]
  wire  acc_io_control_bits_write; // @[AccumulatorWithALUArray.scala 44:19]
  wire  acc_io_tracepoint; // @[AccumulatorWithALUArray.scala 44:19]
  wire [31:0] acc_io_programCounter; // @[AccumulatorWithALUArray.scala 44:19]
  wire  alu_clock; // @[AccumulatorWithALUArray.scala 45:19]
  wire  alu_reset; // @[AccumulatorWithALUArray.scala 45:19]
  wire  alu_io_input_ready; // @[AccumulatorWithALUArray.scala 45:19]
  wire  alu_io_input_valid; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_0; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_1; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_2; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_3; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_4; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_5; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_6; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_7; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_8; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_9; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_10; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_11; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_12; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_13; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_14; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_15; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_16; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_17; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_18; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_19; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_20; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_21; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_22; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_23; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_24; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_25; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_26; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_27; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_28; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_29; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_30; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_input_bits_31; // @[AccumulatorWithALUArray.scala 45:19]
  wire  alu_io_output_ready; // @[AccumulatorWithALUArray.scala 45:19]
  wire  alu_io_output_valid; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_0; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_1; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_2; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_3; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_4; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_5; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_6; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_7; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_8; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_9; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_10; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_11; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_12; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_13; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_14; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_15; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_16; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_17; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_18; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_19; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_20; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_21; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_22; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_23; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_24; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_25; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_26; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_27; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_28; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_29; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_30; // @[AccumulatorWithALUArray.scala 45:19]
  wire [15:0] alu_io_output_bits_31; // @[AccumulatorWithALUArray.scala 45:19]
  wire  alu_io_instruction_ready; // @[AccumulatorWithALUArray.scala 45:19]
  wire  alu_io_instruction_valid; // @[AccumulatorWithALUArray.scala 45:19]
  wire [3:0] alu_io_instruction_bits_op; // @[AccumulatorWithALUArray.scala 45:19]
  wire  alu_io_instruction_bits_sourceLeft; // @[AccumulatorWithALUArray.scala 45:19]
  wire  alu_io_instruction_bits_sourceRight; // @[AccumulatorWithALUArray.scala 45:19]
  wire  alu_io_instruction_bits_dest; // @[AccumulatorWithALUArray.scala 45:19]
  wire  aluOutputDemux_x6_demux_io_in_ready; // @[Demux.scala 46:23]
  wire  aluOutputDemux_x6_demux_io_in_valid; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_0; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_1; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_2; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_3; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_4; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_5; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_6; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_7; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_8; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_9; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_10; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_11; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_12; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_13; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_14; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_15; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_16; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_17; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_18; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_19; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_20; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_21; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_22; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_23; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_24; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_25; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_26; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_27; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_28; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_29; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_30; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_in_bits_31; // @[Demux.scala 46:23]
  wire  aluOutputDemux_x6_demux_io_sel_ready; // @[Demux.scala 46:23]
  wire  aluOutputDemux_x6_demux_io_sel_valid; // @[Demux.scala 46:23]
  wire  aluOutputDemux_x6_demux_io_sel_bits; // @[Demux.scala 46:23]
  wire  aluOutputDemux_x6_demux_io_out_0_ready; // @[Demux.scala 46:23]
  wire  aluOutputDemux_x6_demux_io_out_0_valid; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_0; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_1; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_2; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_3; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_4; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_5; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_6; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_7; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_8; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_9; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_10; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_11; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_12; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_13; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_14; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_15; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_16; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_17; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_18; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_19; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_20; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_21; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_22; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_23; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_24; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_25; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_26; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_27; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_28; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_29; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_30; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_0_bits_31; // @[Demux.scala 46:23]
  wire  aluOutputDemux_x6_demux_io_out_1_ready; // @[Demux.scala 46:23]
  wire  aluOutputDemux_x6_demux_io_out_1_valid; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_0; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_1; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_2; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_3; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_4; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_5; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_6; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_7; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_8; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_9; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_10; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_11; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_12; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_13; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_14; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_15; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_16; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_17; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_18; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_19; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_20; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_21; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_22; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_23; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_24; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_25; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_26; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_27; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_28; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_29; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_30; // @[Demux.scala 46:23]
  wire [15:0] aluOutputDemux_x6_demux_io_out_1_bits_31; // @[Demux.scala 46:23]
  wire  aluOutputDemux_clock; // @[Mem.scala 22:19]
  wire  aluOutputDemux_reset; // @[Mem.scala 22:19]
  wire  aluOutputDemux_io_enq_ready; // @[Mem.scala 22:19]
  wire  aluOutputDemux_io_enq_valid; // @[Mem.scala 22:19]
  wire  aluOutputDemux_io_enq_bits; // @[Mem.scala 22:19]
  wire  aluOutputDemux_io_deq_ready; // @[Mem.scala 22:19]
  wire  aluOutputDemux_io_deq_valid; // @[Mem.scala 22:19]
  wire  aluOutputDemux_io_deq_bits; // @[Mem.scala 22:19]
  wire  accInputMux_x15_mux_io_in_0_ready; // @[Mux.scala 71:21]
  wire  accInputMux_x15_mux_io_in_0_valid; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_0; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_1; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_2; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_3; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_4; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_5; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_6; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_7; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_8; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_9; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_10; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_11; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_12; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_13; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_14; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_15; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_16; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_17; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_18; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_19; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_20; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_21; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_22; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_23; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_24; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_25; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_26; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_27; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_28; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_29; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_30; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_0_bits_31; // @[Mux.scala 71:21]
  wire  accInputMux_x15_mux_io_in_1_ready; // @[Mux.scala 71:21]
  wire  accInputMux_x15_mux_io_in_1_valid; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_0; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_1; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_2; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_3; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_4; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_5; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_6; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_7; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_8; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_9; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_10; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_11; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_12; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_13; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_14; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_15; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_16; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_17; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_18; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_19; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_20; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_21; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_22; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_23; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_24; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_25; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_26; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_27; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_28; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_29; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_30; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_in_1_bits_31; // @[Mux.scala 71:21]
  wire  accInputMux_x15_mux_io_sel_ready; // @[Mux.scala 71:21]
  wire  accInputMux_x15_mux_io_sel_valid; // @[Mux.scala 71:21]
  wire  accInputMux_x15_mux_io_sel_bits; // @[Mux.scala 71:21]
  wire  accInputMux_x15_mux_io_out_ready; // @[Mux.scala 71:21]
  wire  accInputMux_x15_mux_io_out_valid; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_0; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_1; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_2; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_3; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_4; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_5; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_6; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_7; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_8; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_9; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_10; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_11; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_12; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_13; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_14; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_15; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_16; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_17; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_18; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_19; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_20; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_21; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_22; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_23; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_24; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_25; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_26; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_27; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_28; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_29; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_30; // @[Mux.scala 71:21]
  wire [15:0] accInputMux_x15_mux_io_out_bits_31; // @[Mux.scala 71:21]
  wire  accInputMux_clock; // @[Mem.scala 22:19]
  wire  accInputMux_reset; // @[Mem.scala 22:19]
  wire  accInputMux_io_enq_ready; // @[Mem.scala 22:19]
  wire  accInputMux_io_enq_valid; // @[Mem.scala 22:19]
  wire  accInputMux_io_enq_bits; // @[Mem.scala 22:19]
  wire  accInputMux_io_deq_ready; // @[Mem.scala 22:19]
  wire  accInputMux_io_deq_valid; // @[Mem.scala 22:19]
  wire  accInputMux_io_deq_bits; // @[Mem.scala 22:19]
  wire  accOutputDemux_x24_demux_io_in_ready; // @[Demux.scala 46:23]
  wire  accOutputDemux_x24_demux_io_in_valid; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_0; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_1; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_2; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_3; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_4; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_5; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_6; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_7; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_8; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_9; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_10; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_11; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_12; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_13; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_14; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_15; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_16; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_17; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_18; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_19; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_20; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_21; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_22; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_23; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_24; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_25; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_26; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_27; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_28; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_29; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_30; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_in_bits_31; // @[Demux.scala 46:23]
  wire  accOutputDemux_x24_demux_io_sel_ready; // @[Demux.scala 46:23]
  wire  accOutputDemux_x24_demux_io_sel_valid; // @[Demux.scala 46:23]
  wire  accOutputDemux_x24_demux_io_sel_bits; // @[Demux.scala 46:23]
  wire  accOutputDemux_x24_demux_io_out_0_ready; // @[Demux.scala 46:23]
  wire  accOutputDemux_x24_demux_io_out_0_valid; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_0; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_1; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_2; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_3; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_4; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_5; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_6; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_7; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_8; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_9; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_10; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_11; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_12; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_13; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_14; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_15; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_16; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_17; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_18; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_19; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_20; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_21; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_22; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_23; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_24; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_25; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_26; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_27; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_28; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_29; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_30; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_0_bits_31; // @[Demux.scala 46:23]
  wire  accOutputDemux_x24_demux_io_out_1_ready; // @[Demux.scala 46:23]
  wire  accOutputDemux_x24_demux_io_out_1_valid; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_0; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_1; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_2; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_3; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_4; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_5; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_6; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_7; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_8; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_9; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_10; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_11; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_12; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_13; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_14; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_15; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_16; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_17; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_18; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_19; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_20; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_21; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_22; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_23; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_24; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_25; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_26; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_27; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_28; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_29; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_30; // @[Demux.scala 46:23]
  wire [15:0] accOutputDemux_x24_demux_io_out_1_bits_31; // @[Demux.scala 46:23]
  wire  accOutputDemux_clock; // @[Mem.scala 22:19]
  wire  accOutputDemux_reset; // @[Mem.scala 22:19]
  wire  accOutputDemux_io_enq_ready; // @[Mem.scala 22:19]
  wire  accOutputDemux_io_enq_valid; // @[Mem.scala 22:19]
  wire  accOutputDemux_io_enq_bits; // @[Mem.scala 22:19]
  wire  accOutputDemux_io_deq_ready; // @[Mem.scala 22:19]
  wire  accOutputDemux_io_deq_valid; // @[Mem.scala 22:19]
  wire  accOutputDemux_io_deq_bits; // @[Mem.scala 22:19]
  wire  accWriteEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  accWriteEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  accWriteEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  accWriteEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  accWriteEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  accWriteEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  accWriteEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  accWriteEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  accReadEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  accReadEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  accReadEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  accReadEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  accReadEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  accReadEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  accReadEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  accReadEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdRWWriteEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  simdRWWriteEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  simdRWWriteEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdRWWriteEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdRWWriteEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdRWWriteEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdRWWriteEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdRWWriteEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdRWWriteEnqueuer_io_out_2_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdRWWriteEnqueuer_io_out_2_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdRWReadEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  simdRWReadEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  simdRWReadEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdRWReadEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdRWReadEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdRWReadEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdRWReadEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdRWReadEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdRWReadEnqueuer_io_out_2_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdRWReadEnqueuer_io_out_2_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_io_out_2_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_io_out_2_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_io_out_3_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdWriteEnqueuer_io_out_3_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_io_out_2_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_io_out_2_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_io_out_3_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdReadEnqueuer_io_out_3_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  simdEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  simdEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  simdEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  simdEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  reg  readEnqueued; // @[AccumulatorWithALUArray.scala 110:29]
  wire  isNoOp = io_control_bits_instruction_op == 4'h0; // @[AccumulatorWithALUArray.scala 130:44]
  wire  _GEN_10 = readEnqueued & accWriteEnqueuer_io_in_ready; // @[AccumulatorWithALUArray.scala 137:28 138:25 151:25]
  wire  _GEN_26 = io_control_bits_write ? _GEN_10 : accReadEnqueuer_io_in_ready; // @[AccumulatorWithALUArray.scala 136:32 161:23]
  wire  _GEN_42 = io_control_bits_write ? accWriteEnqueuer_io_in_ready : 1'h1; // @[AccumulatorWithALUArray.scala 170:32 171:23 179:23]
  wire  dataPathReady = io_control_bits_read ? _GEN_26 : _GEN_42; // @[AccumulatorWithALUArray.scala 135:29]
  wire  _GEN_0 = dataPathReady ? 1'h0 : readEnqueued; // @[AccumulatorWithALUArray.scala 145:31 146:26 148:26]
  wire  _GEN_1 = readEnqueued & io_control_valid; // @[AccumulatorWithALUArray.scala 137:28 MultiEnqueue.scala 40:17 84:17]
  wire  dataPathReady_acc_io_control_w_ready = acc_io_control_ready; // @[ReadyValid.scala 16:17 MultiEnqueue.scala 85:10]
  wire  _GEN_2 = readEnqueued & dataPathReady_acc_io_control_w_ready; // @[AccumulatorWithALUArray.scala 137:28 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  dataPathReady_acc_io_control_w_valid = accWriteEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  readEnqueued_acc_io_control_w_valid = accReadEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_3 = readEnqueued ? dataPathReady_acc_io_control_w_valid : readEnqueued_acc_io_control_w_valid; // @[AccumulatorWithALUArray.scala 137:28 MultiEnqueue.scala 85:{10,10}]
  wire [11:0] _GEN_4 = readEnqueued ? io_control_bits_writeAddress : io_control_bits_readAddress; // @[AccumulatorWithALUArray.scala 137:28 MultiEnqueue.scala 85:{10,10}]
  wire  _GEN_5 = readEnqueued & io_control_bits_accumulate; // @[AccumulatorWithALUArray.scala 137:28 MultiEnqueue.scala 85:{10,10}]
  wire  dataPathReady_accInputMux_io_enq_w_ready = accInputMux_io_enq_ready; // @[ReadyValid.scala 16:17 MultiEnqueue.scala 86:10]
  wire  _GEN_7 = readEnqueued & dataPathReady_accInputMux_io_enq_w_ready; // @[AccumulatorWithALUArray.scala 137:28 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  dataPathReady_accInputMux_io_enq_w_valid = accWriteEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_8 = readEnqueued & dataPathReady_accInputMux_io_enq_w_valid; // @[AccumulatorWithALUArray.scala 137:28 MultiEnqueue.scala 86:10 package.scala 405:15]
  wire  _GEN_11 = readEnqueued ? _GEN_0 : accReadEnqueuer_io_in_ready; // @[AccumulatorWithALUArray.scala 137:28 152:24]
  wire  _GEN_12 = readEnqueued ? 1'h0 : io_control_valid; // @[AccumulatorWithALUArray.scala 137:28 MultiEnqueue.scala 40:17 84:17]
  wire  _GEN_13 = readEnqueued ? 1'h0 : dataPathReady_acc_io_control_w_ready; // @[AccumulatorWithALUArray.scala 137:28 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  readEnqueued_accOutputDemux_io_enq_w_ready = accOutputDemux_io_enq_ready; // @[ReadyValid.scala 16:17 MultiEnqueue.scala 86:10]
  wire  _GEN_14 = readEnqueued ? 1'h0 : readEnqueued_accOutputDemux_io_enq_w_ready; // @[AccumulatorWithALUArray.scala 137:28 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  readEnqueued_accOutputDemux_io_enq_w_valid = accReadEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_15 = readEnqueued ? 1'h0 : readEnqueued_accOutputDemux_io_enq_w_valid; // @[AccumulatorWithALUArray.scala 137:28 package.scala 405:15 MultiEnqueue.scala 86:10]
  wire  _GEN_17 = io_control_bits_write & _GEN_1; // @[AccumulatorWithALUArray.scala 136:32 MultiEnqueue.scala 40:17]
  wire  _GEN_18 = io_control_bits_write & _GEN_2; // @[AccumulatorWithALUArray.scala 136:32 MultiEnqueue.scala 42:18]
  wire  _GEN_19 = io_control_bits_write ? _GEN_3 : readEnqueued_acc_io_control_w_valid; // @[AccumulatorWithALUArray.scala 136:32 MultiEnqueue.scala 85:10]
  wire [11:0] _GEN_20 = io_control_bits_write ? _GEN_4 : io_control_bits_readAddress; // @[AccumulatorWithALUArray.scala 136:32 MultiEnqueue.scala 85:10]
  wire  _GEN_21 = io_control_bits_write & _GEN_5; // @[AccumulatorWithALUArray.scala 136:32 MultiEnqueue.scala 85:10]
  wire  _GEN_22 = io_control_bits_write & readEnqueued; // @[AccumulatorWithALUArray.scala 136:32 MultiEnqueue.scala 85:10]
  wire  _GEN_23 = io_control_bits_write & _GEN_7; // @[AccumulatorWithALUArray.scala 136:32 MultiEnqueue.scala 42:18]
  wire  _GEN_24 = io_control_bits_write & _GEN_8; // @[AccumulatorWithALUArray.scala 136:32 package.scala 405:15]
  wire  _GEN_27 = io_control_bits_write & _GEN_11; // @[AccumulatorWithALUArray.scala 111:16 136:32]
  wire  _GEN_28 = io_control_bits_write ? _GEN_12 : io_control_valid; // @[AccumulatorWithALUArray.scala 136:32 MultiEnqueue.scala 84:17]
  wire  _GEN_29 = io_control_bits_write ? _GEN_13 : dataPathReady_acc_io_control_w_ready; // @[AccumulatorWithALUArray.scala 136:32 ReadyValid.scala 19:11]
  wire  _GEN_30 = io_control_bits_write ? _GEN_14 : readEnqueued_accOutputDemux_io_enq_w_ready; // @[AccumulatorWithALUArray.scala 136:32 ReadyValid.scala 19:11]
  wire  _GEN_31 = io_control_bits_write ? _GEN_15 : readEnqueued_accOutputDemux_io_enq_w_valid; // @[AccumulatorWithALUArray.scala 136:32 MultiEnqueue.scala 86:10]
  wire  _GEN_33 = io_control_bits_write & io_control_valid; // @[AccumulatorWithALUArray.scala 170:32 MultiEnqueue.scala 40:17 84:17]
  wire  _GEN_34 = io_control_bits_write & dataPathReady_acc_io_control_w_ready; // @[AccumulatorWithALUArray.scala 170:32 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  _GEN_35 = io_control_bits_write & dataPathReady_acc_io_control_w_valid; // @[AccumulatorWithALUArray.scala 170:32 MultiEnqueue.scala 85:10 package.scala 405:15]
  wire [11:0] _GEN_36 = io_control_bits_write ? io_control_bits_writeAddress : 12'h0; // @[AccumulatorWithALUArray.scala 170:32 MultiEnqueue.scala 85:10 package.scala 404:14]
  wire  _GEN_37 = io_control_bits_write & io_control_bits_accumulate; // @[AccumulatorWithALUArray.scala 170:32 MultiEnqueue.scala 85:10 package.scala 404:14]
  wire  _GEN_39 = io_control_bits_write & dataPathReady_accInputMux_io_enq_w_ready; // @[AccumulatorWithALUArray.scala 170:32 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  _GEN_40 = io_control_bits_write & dataPathReady_accInputMux_io_enq_w_valid; // @[AccumulatorWithALUArray.scala 170:32 MultiEnqueue.scala 86:10 package.scala 405:15]
  wire  _GEN_43 = io_control_bits_read ? _GEN_17 : _GEN_33; // @[AccumulatorWithALUArray.scala 135:29]
  wire  _GEN_44 = io_control_bits_read ? _GEN_18 : _GEN_34; // @[AccumulatorWithALUArray.scala 135:29]
  wire  _GEN_45 = io_control_bits_read ? _GEN_19 : _GEN_35; // @[AccumulatorWithALUArray.scala 135:29]
  wire [11:0] _GEN_46 = io_control_bits_read ? _GEN_20 : _GEN_36; // @[AccumulatorWithALUArray.scala 135:29]
  wire  _GEN_47 = io_control_bits_read ? _GEN_21 : _GEN_37; // @[AccumulatorWithALUArray.scala 135:29]
  wire  _GEN_48 = io_control_bits_read ? _GEN_22 : io_control_bits_write; // @[AccumulatorWithALUArray.scala 135:29]
  wire  _GEN_49 = io_control_bits_read ? _GEN_23 : _GEN_39; // @[AccumulatorWithALUArray.scala 135:29]
  wire  _GEN_50 = io_control_bits_read ? _GEN_24 : _GEN_40; // @[AccumulatorWithALUArray.scala 135:29]
  wire  _GEN_53 = io_control_bits_read & _GEN_27; // @[AccumulatorWithALUArray.scala 111:16 135:29]
  wire  _GEN_54 = io_control_bits_read & _GEN_28; // @[AccumulatorWithALUArray.scala 135:29 MultiEnqueue.scala 40:17]
  wire  _GEN_55 = io_control_bits_read & _GEN_29; // @[AccumulatorWithALUArray.scala 135:29 MultiEnqueue.scala 42:18]
  wire  _GEN_56 = io_control_bits_read & _GEN_30; // @[AccumulatorWithALUArray.scala 135:29 MultiEnqueue.scala 42:18]
  wire  _GEN_57 = io_control_bits_read & _GEN_31; // @[AccumulatorWithALUArray.scala 135:29 package.scala 405:15]
  wire  _GEN_87 = readEnqueued & simdRWWriteEnqueuer_io_in_ready; // @[AccumulatorWithALUArray.scala 188:28 189:25 204:25]
  wire  _GEN_111 = io_control_bits_write ? _GEN_87 : simdReadEnqueuer_io_in_ready; // @[AccumulatorWithALUArray.scala 186:32 222:23]
  wire  _GEN_146 = io_control_bits_write ? simdWriteEnqueuer_io_in_ready : simdEnqueuer_io_in_ready; // @[AccumulatorWithALUArray.scala 235:32 236:23 248:23]
  wire  dataPathReady_1 = io_control_bits_read ? _GEN_111 : _GEN_146; // @[AccumulatorWithALUArray.scala 185:29]
  wire  _GEN_59 = dataPathReady_1 ? 1'h0 : readEnqueued; // @[AccumulatorWithALUArray.scala 198:31 199:26 201:26]
  wire  _T_2 = ~io_control_bits_instruction_sourceLeft | ~io_control_bits_instruction_sourceRight; // @[AccumulatorWithALUArray.scala 206:57]
  wire  _GEN_60 = _T_2 & io_control_valid; // @[AccumulatorWithALUArray.scala 207:13 MultiEnqueue.scala 114:17 40:17]
  wire  _GEN_61 = _T_2 & dataPathReady_acc_io_control_w_ready; // @[AccumulatorWithALUArray.scala 207:13 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  readEnqueued_acc_io_control_w_1_valid = simdRWReadEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_62 = _T_2 & readEnqueued_acc_io_control_w_1_valid; // @[AccumulatorWithALUArray.scala 207:13 MultiEnqueue.scala 115:10 package.scala 405:15]
  wire [11:0] _GEN_63 = _T_2 ? io_control_bits_readAddress : 12'h0; // @[AccumulatorWithALUArray.scala 207:13 MultiEnqueue.scala 115:10 package.scala 404:14]
  wire  _GEN_66 = _T_2 & readEnqueued_accOutputDemux_io_enq_w_ready; // @[AccumulatorWithALUArray.scala 207:13 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  readEnqueued_accOutputDemux_io_enq_w_1_valid = simdRWReadEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_67 = _T_2 & readEnqueued_accOutputDemux_io_enq_w_1_valid; // @[AccumulatorWithALUArray.scala 207:13 MultiEnqueue.scala 116:10 package.scala 405:15]
  wire  readEnqueued_alu_io_instruction_w_ready = alu_io_instruction_ready; // @[MultiEnqueue.scala 117:10 ReadyValid.scala 16:17]
  wire  _GEN_69 = _T_2 & readEnqueued_alu_io_instruction_w_ready; // @[AccumulatorWithALUArray.scala 207:13 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  readEnqueued_alu_io_instruction_w_valid = simdRWReadEnqueuer_io_out_2_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_70 = _T_2 & readEnqueued_alu_io_instruction_w_valid; // @[AccumulatorWithALUArray.scala 207:13 MultiEnqueue.scala 117:10 package.scala 405:15]
  wire [3:0] _GEN_71 = _T_2 ? io_control_bits_instruction_op : 4'h0; // @[AccumulatorWithALUArray.scala 207:13 MultiEnqueue.scala 117:10 package.scala 404:14]
  wire  _GEN_72 = _T_2 & io_control_bits_instruction_sourceLeft; // @[AccumulatorWithALUArray.scala 207:13 MultiEnqueue.scala 117:10 package.scala 404:14]
  wire  _GEN_73 = _T_2 & io_control_bits_instruction_sourceRight; // @[AccumulatorWithALUArray.scala 207:13 MultiEnqueue.scala 117:10 package.scala 404:14]
  wire  _GEN_74 = _T_2 & io_control_bits_instruction_dest; // @[AccumulatorWithALUArray.scala 207:13 MultiEnqueue.scala 117:10 package.scala 404:14]
  wire  _GEN_75 = _T_2 ? simdRWReadEnqueuer_io_in_ready : 1'h1; // @[AccumulatorWithALUArray.scala 207:13 208:26 218:26]
  wire  dataPathReady_acc_io_control_w_3_valid = simdRWWriteEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_77 = readEnqueued ? dataPathReady_acc_io_control_w_3_valid : _GEN_62; // @[AccumulatorWithALUArray.scala 188:28 MultiEnqueue.scala 115:10]
  wire [11:0] _GEN_78 = readEnqueued ? io_control_bits_writeAddress : _GEN_63; // @[AccumulatorWithALUArray.scala 188:28 MultiEnqueue.scala 115:10]
  wire  dataPathReady_aluOutputDemux_io_enq_w_ready = aluOutputDemux_io_enq_ready; // @[MultiEnqueue.scala 116:10 ReadyValid.scala 16:17]
  wire  _GEN_81 = readEnqueued & dataPathReady_aluOutputDemux_io_enq_w_ready; // @[AccumulatorWithALUArray.scala 188:28 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  dataPathReady_aluOutputDemux_io_enq_w_valid = simdRWWriteEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_82 = readEnqueued & dataPathReady_aluOutputDemux_io_enq_w_valid; // @[AccumulatorWithALUArray.scala 188:28 MultiEnqueue.scala 116:10 package.scala 405:15]
  wire  dataPathReady_accInputMux_io_enq_w_2_valid = simdRWWriteEnqueuer_io_out_2_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_85 = readEnqueued & dataPathReady_accInputMux_io_enq_w_2_valid; // @[AccumulatorWithALUArray.scala 188:28 MultiEnqueue.scala 117:10 package.scala 405:15]
  wire  _GEN_88 = readEnqueued ? _GEN_59 : _GEN_75; // @[AccumulatorWithALUArray.scala 188:28]
  wire  _GEN_89 = readEnqueued ? 1'h0 : _GEN_60; // @[AccumulatorWithALUArray.scala 188:28 MultiEnqueue.scala 40:17]
  wire  _GEN_90 = readEnqueued ? 1'h0 : _GEN_61; // @[AccumulatorWithALUArray.scala 188:28 MultiEnqueue.scala 42:18]
  wire  _GEN_91 = readEnqueued ? 1'h0 : _GEN_66; // @[AccumulatorWithALUArray.scala 188:28 MultiEnqueue.scala 42:18]
  wire  _GEN_92 = readEnqueued ? 1'h0 : _GEN_67; // @[AccumulatorWithALUArray.scala 188:28 package.scala 405:15]
  wire  _GEN_93 = readEnqueued ? 1'h0 : _T_2; // @[AccumulatorWithALUArray.scala 188:28 package.scala 404:14]
  wire  _GEN_94 = readEnqueued ? 1'h0 : _GEN_69; // @[AccumulatorWithALUArray.scala 188:28 MultiEnqueue.scala 42:18]
  wire  _GEN_95 = readEnqueued ? 1'h0 : _GEN_70; // @[AccumulatorWithALUArray.scala 188:28 package.scala 405:15]
  wire [3:0] _GEN_96 = readEnqueued ? 4'h0 : _GEN_71; // @[AccumulatorWithALUArray.scala 188:28 package.scala 404:14]
  wire  _GEN_97 = readEnqueued ? 1'h0 : _GEN_72; // @[AccumulatorWithALUArray.scala 188:28 package.scala 404:14]
  wire  _GEN_98 = readEnqueued ? 1'h0 : _GEN_73; // @[AccumulatorWithALUArray.scala 188:28 package.scala 404:14]
  wire  _GEN_99 = readEnqueued ? 1'h0 : _GEN_74; // @[AccumulatorWithALUArray.scala 188:28 package.scala 404:14]
  wire  dataPathReady_acc_io_control_w_4_valid = simdReadEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_101 = io_control_bits_write ? _GEN_77 : dataPathReady_acc_io_control_w_4_valid; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 151:10]
  wire [11:0] _GEN_102 = io_control_bits_write ? _GEN_78 : io_control_bits_readAddress; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 151:10]
  wire  _GEN_105 = io_control_bits_write & _GEN_81; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 42:18]
  wire  dataPathReady_aluOutputDemux_io_enq_w_1_valid = simdReadEnqueuer_io_out_2_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_106 = io_control_bits_write ? _GEN_82 : dataPathReady_aluOutputDemux_io_enq_w_1_valid; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 153:10]
  wire  _GEN_109 = io_control_bits_write & _GEN_85; // @[AccumulatorWithALUArray.scala 186:32 package.scala 405:15]
  wire  _GEN_112 = io_control_bits_write & _GEN_88; // @[AccumulatorWithALUArray.scala 111:16 186:32]
  wire  _GEN_113 = io_control_bits_write & _GEN_89; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 40:17]
  wire  _GEN_114 = io_control_bits_write & _GEN_90; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 42:18]
  wire  _GEN_115 = io_control_bits_write & _GEN_91; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 42:18]
  wire  dataPathReady_accOutputDemux_io_enq_w_1_valid = simdReadEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_116 = io_control_bits_write ? _GEN_92 : dataPathReady_accOutputDemux_io_enq_w_1_valid; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 152:10]
  wire  _GEN_117 = io_control_bits_write ? _GEN_93 : 1'h1; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 152:10]
  wire  _GEN_118 = io_control_bits_write & _GEN_94; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 42:18]
  wire  dataPathReady_alu_io_instruction_w_valid = simdReadEnqueuer_io_out_3_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_119 = io_control_bits_write ? _GEN_95 : dataPathReady_alu_io_instruction_w_valid; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 154:10]
  wire [3:0] _GEN_120 = io_control_bits_write ? _GEN_96 : io_control_bits_instruction_op; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 154:10]
  wire  _GEN_121 = io_control_bits_write ? _GEN_97 : io_control_bits_instruction_sourceLeft; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 154:10]
  wire  _GEN_122 = io_control_bits_write ? _GEN_98 : io_control_bits_instruction_sourceRight; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 154:10]
  wire  _GEN_123 = io_control_bits_write ? _GEN_99 : io_control_bits_instruction_dest; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 154:10]
  wire  _GEN_124 = io_control_bits_write ? 1'h0 : io_control_valid; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 150:17 40:17]
  wire  _GEN_125 = io_control_bits_write ? 1'h0 : dataPathReady_acc_io_control_w_ready; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  _GEN_126 = io_control_bits_write ? 1'h0 : readEnqueued_accOutputDemux_io_enq_w_ready; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  _GEN_127 = io_control_bits_write ? 1'h0 : dataPathReady_aluOutputDemux_io_enq_w_ready; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  _GEN_128 = io_control_bits_write ? 1'h0 : readEnqueued_alu_io_instruction_w_ready; // @[AccumulatorWithALUArray.scala 186:32 MultiEnqueue.scala 42:18 ReadyValid.scala 19:11]
  wire  dataPathReady_acc_io_control_w_5_valid = simdWriteEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_130 = io_control_bits_write & dataPathReady_acc_io_control_w_5_valid; // @[AccumulatorWithALUArray.scala 235:32 MultiEnqueue.scala 151:10 package.scala 405:15]
  wire  _GEN_134 = io_control_bits_write & dataPathReady_aluOutputDemux_io_enq_w_ready; // @[AccumulatorWithALUArray.scala 235:32 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  dataPathReady_aluOutputDemux_io_enq_w_2_valid = simdWriteEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  dataPathReady_aluOutputDemux_io_enq_w_3_valid = simdEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_135 = io_control_bits_write ? dataPathReady_aluOutputDemux_io_enq_w_2_valid :
    dataPathReady_aluOutputDemux_io_enq_w_3_valid; // @[AccumulatorWithALUArray.scala 235:32 MultiEnqueue.scala 152:10 85:10]
  wire  dataPathReady_accInputMux_io_enq_w_3_valid = simdWriteEnqueuer_io_out_2_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_138 = io_control_bits_write & dataPathReady_accInputMux_io_enq_w_3_valid; // @[AccumulatorWithALUArray.scala 235:32 MultiEnqueue.scala 153:10 package.scala 405:15]
  wire  _GEN_140 = io_control_bits_write & readEnqueued_alu_io_instruction_w_ready; // @[AccumulatorWithALUArray.scala 235:32 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  dataPathReady_alu_io_instruction_w_1_valid = simdWriteEnqueuer_io_out_3_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  dataPathReady_alu_io_instruction_w_2_valid = simdEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_141 = io_control_bits_write ? dataPathReady_alu_io_instruction_w_1_valid :
    dataPathReady_alu_io_instruction_w_2_valid; // @[AccumulatorWithALUArray.scala 235:32 MultiEnqueue.scala 154:10 86:10]
  wire  _GEN_149 = io_control_bits_read & _GEN_17; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 40:17]
  wire  _GEN_150 = io_control_bits_read & _GEN_18; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_151 = io_control_bits_read ? _GEN_101 : _GEN_130; // @[AccumulatorWithALUArray.scala 185:29]
  wire [11:0] _GEN_152 = io_control_bits_read ? _GEN_102 : _GEN_36; // @[AccumulatorWithALUArray.scala 185:29]
  wire  _GEN_155 = io_control_bits_read & _GEN_105; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_156 = io_control_bits_read ? _GEN_106 : _GEN_135; // @[AccumulatorWithALUArray.scala 185:29]
  wire  _GEN_158 = io_control_bits_read & _GEN_23; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_159 = io_control_bits_read ? _GEN_109 : _GEN_138; // @[AccumulatorWithALUArray.scala 185:29]
  wire  _GEN_162 = io_control_bits_read & _GEN_112; // @[AccumulatorWithALUArray.scala 111:16 185:29]
  wire  _GEN_163 = io_control_bits_read & _GEN_113; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 40:17]
  wire  _GEN_164 = io_control_bits_read & _GEN_114; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_165 = io_control_bits_read & _GEN_115; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_166 = io_control_bits_read & _GEN_116; // @[AccumulatorWithALUArray.scala 185:29 package.scala 405:15]
  wire  _GEN_167 = io_control_bits_read & _GEN_117; // @[AccumulatorWithALUArray.scala 185:29 package.scala 404:14]
  wire  _GEN_168 = io_control_bits_read & _GEN_118; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_169 = io_control_bits_read ? _GEN_119 : _GEN_141; // @[AccumulatorWithALUArray.scala 185:29]
  wire [3:0] _GEN_170 = io_control_bits_read ? _GEN_120 : io_control_bits_instruction_op; // @[AccumulatorWithALUArray.scala 185:29]
  wire  _GEN_171 = io_control_bits_read ? _GEN_121 : io_control_bits_instruction_sourceLeft; // @[AccumulatorWithALUArray.scala 185:29]
  wire  _GEN_172 = io_control_bits_read ? _GEN_122 : io_control_bits_instruction_sourceRight; // @[AccumulatorWithALUArray.scala 185:29]
  wire  _GEN_173 = io_control_bits_read ? _GEN_123 : io_control_bits_instruction_dest; // @[AccumulatorWithALUArray.scala 185:29]
  wire  _GEN_174 = io_control_bits_read & _GEN_124; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 40:17]
  wire  _GEN_175 = io_control_bits_read & _GEN_125; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_176 = io_control_bits_read & _GEN_126; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_177 = io_control_bits_read & _GEN_127; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_178 = io_control_bits_read & _GEN_128; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_179 = io_control_bits_read ? 1'h0 : _GEN_33; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 40:17]
  wire  _GEN_180 = io_control_bits_read ? 1'h0 : _GEN_34; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_181 = io_control_bits_read ? 1'h0 : _GEN_134; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_182 = io_control_bits_read ? 1'h0 : _GEN_39; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_183 = io_control_bits_read ? 1'h0 : _GEN_140; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_184 = io_control_bits_read ? 1'h0 : _GEN_124; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 40:17]
  wire  _GEN_185 = io_control_bits_read ? 1'h0 : _GEN_127; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  wire  _GEN_186 = io_control_bits_read ? 1'h0 : _GEN_128; // @[AccumulatorWithALUArray.scala 185:29 MultiEnqueue.scala 42:18]
  Accumulator acc ( // @[AccumulatorWithALUArray.scala 44:19]
    .clock(acc_clock),
    .reset(acc_reset),
    .io_input_ready(acc_io_input_ready),
    .io_input_valid(acc_io_input_valid),
    .io_input_bits_0(acc_io_input_bits_0),
    .io_input_bits_1(acc_io_input_bits_1),
    .io_input_bits_2(acc_io_input_bits_2),
    .io_input_bits_3(acc_io_input_bits_3),
    .io_input_bits_4(acc_io_input_bits_4),
    .io_input_bits_5(acc_io_input_bits_5),
    .io_input_bits_6(acc_io_input_bits_6),
    .io_input_bits_7(acc_io_input_bits_7),
    .io_input_bits_8(acc_io_input_bits_8),
    .io_input_bits_9(acc_io_input_bits_9),
    .io_input_bits_10(acc_io_input_bits_10),
    .io_input_bits_11(acc_io_input_bits_11),
    .io_input_bits_12(acc_io_input_bits_12),
    .io_input_bits_13(acc_io_input_bits_13),
    .io_input_bits_14(acc_io_input_bits_14),
    .io_input_bits_15(acc_io_input_bits_15),
    .io_input_bits_16(acc_io_input_bits_16),
    .io_input_bits_17(acc_io_input_bits_17),
    .io_input_bits_18(acc_io_input_bits_18),
    .io_input_bits_19(acc_io_input_bits_19),
    .io_input_bits_20(acc_io_input_bits_20),
    .io_input_bits_21(acc_io_input_bits_21),
    .io_input_bits_22(acc_io_input_bits_22),
    .io_input_bits_23(acc_io_input_bits_23),
    .io_input_bits_24(acc_io_input_bits_24),
    .io_input_bits_25(acc_io_input_bits_25),
    .io_input_bits_26(acc_io_input_bits_26),
    .io_input_bits_27(acc_io_input_bits_27),
    .io_input_bits_28(acc_io_input_bits_28),
    .io_input_bits_29(acc_io_input_bits_29),
    .io_input_bits_30(acc_io_input_bits_30),
    .io_input_bits_31(acc_io_input_bits_31),
    .io_output_ready(acc_io_output_ready),
    .io_output_valid(acc_io_output_valid),
    .io_output_bits_0(acc_io_output_bits_0),
    .io_output_bits_1(acc_io_output_bits_1),
    .io_output_bits_2(acc_io_output_bits_2),
    .io_output_bits_3(acc_io_output_bits_3),
    .io_output_bits_4(acc_io_output_bits_4),
    .io_output_bits_5(acc_io_output_bits_5),
    .io_output_bits_6(acc_io_output_bits_6),
    .io_output_bits_7(acc_io_output_bits_7),
    .io_output_bits_8(acc_io_output_bits_8),
    .io_output_bits_9(acc_io_output_bits_9),
    .io_output_bits_10(acc_io_output_bits_10),
    .io_output_bits_11(acc_io_output_bits_11),
    .io_output_bits_12(acc_io_output_bits_12),
    .io_output_bits_13(acc_io_output_bits_13),
    .io_output_bits_14(acc_io_output_bits_14),
    .io_output_bits_15(acc_io_output_bits_15),
    .io_output_bits_16(acc_io_output_bits_16),
    .io_output_bits_17(acc_io_output_bits_17),
    .io_output_bits_18(acc_io_output_bits_18),
    .io_output_bits_19(acc_io_output_bits_19),
    .io_output_bits_20(acc_io_output_bits_20),
    .io_output_bits_21(acc_io_output_bits_21),
    .io_output_bits_22(acc_io_output_bits_22),
    .io_output_bits_23(acc_io_output_bits_23),
    .io_output_bits_24(acc_io_output_bits_24),
    .io_output_bits_25(acc_io_output_bits_25),
    .io_output_bits_26(acc_io_output_bits_26),
    .io_output_bits_27(acc_io_output_bits_27),
    .io_output_bits_28(acc_io_output_bits_28),
    .io_output_bits_29(acc_io_output_bits_29),
    .io_output_bits_30(acc_io_output_bits_30),
    .io_output_bits_31(acc_io_output_bits_31),
    .io_control_ready(acc_io_control_ready),
    .io_control_valid(acc_io_control_valid),
    .io_control_bits_address(acc_io_control_bits_address),
    .io_control_bits_accumulate(acc_io_control_bits_accumulate),
    .io_control_bits_write(acc_io_control_bits_write),
    .io_tracepoint(acc_io_tracepoint),
    .io_programCounter(acc_io_programCounter)
  );
  ALUArray alu ( // @[AccumulatorWithALUArray.scala 45:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_input_ready(alu_io_input_ready),
    .io_input_valid(alu_io_input_valid),
    .io_input_bits_0(alu_io_input_bits_0),
    .io_input_bits_1(alu_io_input_bits_1),
    .io_input_bits_2(alu_io_input_bits_2),
    .io_input_bits_3(alu_io_input_bits_3),
    .io_input_bits_4(alu_io_input_bits_4),
    .io_input_bits_5(alu_io_input_bits_5),
    .io_input_bits_6(alu_io_input_bits_6),
    .io_input_bits_7(alu_io_input_bits_7),
    .io_input_bits_8(alu_io_input_bits_8),
    .io_input_bits_9(alu_io_input_bits_9),
    .io_input_bits_10(alu_io_input_bits_10),
    .io_input_bits_11(alu_io_input_bits_11),
    .io_input_bits_12(alu_io_input_bits_12),
    .io_input_bits_13(alu_io_input_bits_13),
    .io_input_bits_14(alu_io_input_bits_14),
    .io_input_bits_15(alu_io_input_bits_15),
    .io_input_bits_16(alu_io_input_bits_16),
    .io_input_bits_17(alu_io_input_bits_17),
    .io_input_bits_18(alu_io_input_bits_18),
    .io_input_bits_19(alu_io_input_bits_19),
    .io_input_bits_20(alu_io_input_bits_20),
    .io_input_bits_21(alu_io_input_bits_21),
    .io_input_bits_22(alu_io_input_bits_22),
    .io_input_bits_23(alu_io_input_bits_23),
    .io_input_bits_24(alu_io_input_bits_24),
    .io_input_bits_25(alu_io_input_bits_25),
    .io_input_bits_26(alu_io_input_bits_26),
    .io_input_bits_27(alu_io_input_bits_27),
    .io_input_bits_28(alu_io_input_bits_28),
    .io_input_bits_29(alu_io_input_bits_29),
    .io_input_bits_30(alu_io_input_bits_30),
    .io_input_bits_31(alu_io_input_bits_31),
    .io_output_ready(alu_io_output_ready),
    .io_output_valid(alu_io_output_valid),
    .io_output_bits_0(alu_io_output_bits_0),
    .io_output_bits_1(alu_io_output_bits_1),
    .io_output_bits_2(alu_io_output_bits_2),
    .io_output_bits_3(alu_io_output_bits_3),
    .io_output_bits_4(alu_io_output_bits_4),
    .io_output_bits_5(alu_io_output_bits_5),
    .io_output_bits_6(alu_io_output_bits_6),
    .io_output_bits_7(alu_io_output_bits_7),
    .io_output_bits_8(alu_io_output_bits_8),
    .io_output_bits_9(alu_io_output_bits_9),
    .io_output_bits_10(alu_io_output_bits_10),
    .io_output_bits_11(alu_io_output_bits_11),
    .io_output_bits_12(alu_io_output_bits_12),
    .io_output_bits_13(alu_io_output_bits_13),
    .io_output_bits_14(alu_io_output_bits_14),
    .io_output_bits_15(alu_io_output_bits_15),
    .io_output_bits_16(alu_io_output_bits_16),
    .io_output_bits_17(alu_io_output_bits_17),
    .io_output_bits_18(alu_io_output_bits_18),
    .io_output_bits_19(alu_io_output_bits_19),
    .io_output_bits_20(alu_io_output_bits_20),
    .io_output_bits_21(alu_io_output_bits_21),
    .io_output_bits_22(alu_io_output_bits_22),
    .io_output_bits_23(alu_io_output_bits_23),
    .io_output_bits_24(alu_io_output_bits_24),
    .io_output_bits_25(alu_io_output_bits_25),
    .io_output_bits_26(alu_io_output_bits_26),
    .io_output_bits_27(alu_io_output_bits_27),
    .io_output_bits_28(alu_io_output_bits_28),
    .io_output_bits_29(alu_io_output_bits_29),
    .io_output_bits_30(alu_io_output_bits_30),
    .io_output_bits_31(alu_io_output_bits_31),
    .io_instruction_ready(alu_io_instruction_ready),
    .io_instruction_valid(alu_io_instruction_valid),
    .io_instruction_bits_op(alu_io_instruction_bits_op),
    .io_instruction_bits_sourceLeft(alu_io_instruction_bits_sourceLeft),
    .io_instruction_bits_sourceRight(alu_io_instruction_bits_sourceRight),
    .io_instruction_bits_dest(alu_io_instruction_bits_dest)
  );
  Demux aluOutputDemux_x6_demux ( // @[Demux.scala 46:23]
    .io_in_ready(aluOutputDemux_x6_demux_io_in_ready),
    .io_in_valid(aluOutputDemux_x6_demux_io_in_valid),
    .io_in_bits_0(aluOutputDemux_x6_demux_io_in_bits_0),
    .io_in_bits_1(aluOutputDemux_x6_demux_io_in_bits_1),
    .io_in_bits_2(aluOutputDemux_x6_demux_io_in_bits_2),
    .io_in_bits_3(aluOutputDemux_x6_demux_io_in_bits_3),
    .io_in_bits_4(aluOutputDemux_x6_demux_io_in_bits_4),
    .io_in_bits_5(aluOutputDemux_x6_demux_io_in_bits_5),
    .io_in_bits_6(aluOutputDemux_x6_demux_io_in_bits_6),
    .io_in_bits_7(aluOutputDemux_x6_demux_io_in_bits_7),
    .io_in_bits_8(aluOutputDemux_x6_demux_io_in_bits_8),
    .io_in_bits_9(aluOutputDemux_x6_demux_io_in_bits_9),
    .io_in_bits_10(aluOutputDemux_x6_demux_io_in_bits_10),
    .io_in_bits_11(aluOutputDemux_x6_demux_io_in_bits_11),
    .io_in_bits_12(aluOutputDemux_x6_demux_io_in_bits_12),
    .io_in_bits_13(aluOutputDemux_x6_demux_io_in_bits_13),
    .io_in_bits_14(aluOutputDemux_x6_demux_io_in_bits_14),
    .io_in_bits_15(aluOutputDemux_x6_demux_io_in_bits_15),
    .io_in_bits_16(aluOutputDemux_x6_demux_io_in_bits_16),
    .io_in_bits_17(aluOutputDemux_x6_demux_io_in_bits_17),
    .io_in_bits_18(aluOutputDemux_x6_demux_io_in_bits_18),
    .io_in_bits_19(aluOutputDemux_x6_demux_io_in_bits_19),
    .io_in_bits_20(aluOutputDemux_x6_demux_io_in_bits_20),
    .io_in_bits_21(aluOutputDemux_x6_demux_io_in_bits_21),
    .io_in_bits_22(aluOutputDemux_x6_demux_io_in_bits_22),
    .io_in_bits_23(aluOutputDemux_x6_demux_io_in_bits_23),
    .io_in_bits_24(aluOutputDemux_x6_demux_io_in_bits_24),
    .io_in_bits_25(aluOutputDemux_x6_demux_io_in_bits_25),
    .io_in_bits_26(aluOutputDemux_x6_demux_io_in_bits_26),
    .io_in_bits_27(aluOutputDemux_x6_demux_io_in_bits_27),
    .io_in_bits_28(aluOutputDemux_x6_demux_io_in_bits_28),
    .io_in_bits_29(aluOutputDemux_x6_demux_io_in_bits_29),
    .io_in_bits_30(aluOutputDemux_x6_demux_io_in_bits_30),
    .io_in_bits_31(aluOutputDemux_x6_demux_io_in_bits_31),
    .io_sel_ready(aluOutputDemux_x6_demux_io_sel_ready),
    .io_sel_valid(aluOutputDemux_x6_demux_io_sel_valid),
    .io_sel_bits(aluOutputDemux_x6_demux_io_sel_bits),
    .io_out_0_ready(aluOutputDemux_x6_demux_io_out_0_ready),
    .io_out_0_valid(aluOutputDemux_x6_demux_io_out_0_valid),
    .io_out_0_bits_0(aluOutputDemux_x6_demux_io_out_0_bits_0),
    .io_out_0_bits_1(aluOutputDemux_x6_demux_io_out_0_bits_1),
    .io_out_0_bits_2(aluOutputDemux_x6_demux_io_out_0_bits_2),
    .io_out_0_bits_3(aluOutputDemux_x6_demux_io_out_0_bits_3),
    .io_out_0_bits_4(aluOutputDemux_x6_demux_io_out_0_bits_4),
    .io_out_0_bits_5(aluOutputDemux_x6_demux_io_out_0_bits_5),
    .io_out_0_bits_6(aluOutputDemux_x6_demux_io_out_0_bits_6),
    .io_out_0_bits_7(aluOutputDemux_x6_demux_io_out_0_bits_7),
    .io_out_0_bits_8(aluOutputDemux_x6_demux_io_out_0_bits_8),
    .io_out_0_bits_9(aluOutputDemux_x6_demux_io_out_0_bits_9),
    .io_out_0_bits_10(aluOutputDemux_x6_demux_io_out_0_bits_10),
    .io_out_0_bits_11(aluOutputDemux_x6_demux_io_out_0_bits_11),
    .io_out_0_bits_12(aluOutputDemux_x6_demux_io_out_0_bits_12),
    .io_out_0_bits_13(aluOutputDemux_x6_demux_io_out_0_bits_13),
    .io_out_0_bits_14(aluOutputDemux_x6_demux_io_out_0_bits_14),
    .io_out_0_bits_15(aluOutputDemux_x6_demux_io_out_0_bits_15),
    .io_out_0_bits_16(aluOutputDemux_x6_demux_io_out_0_bits_16),
    .io_out_0_bits_17(aluOutputDemux_x6_demux_io_out_0_bits_17),
    .io_out_0_bits_18(aluOutputDemux_x6_demux_io_out_0_bits_18),
    .io_out_0_bits_19(aluOutputDemux_x6_demux_io_out_0_bits_19),
    .io_out_0_bits_20(aluOutputDemux_x6_demux_io_out_0_bits_20),
    .io_out_0_bits_21(aluOutputDemux_x6_demux_io_out_0_bits_21),
    .io_out_0_bits_22(aluOutputDemux_x6_demux_io_out_0_bits_22),
    .io_out_0_bits_23(aluOutputDemux_x6_demux_io_out_0_bits_23),
    .io_out_0_bits_24(aluOutputDemux_x6_demux_io_out_0_bits_24),
    .io_out_0_bits_25(aluOutputDemux_x6_demux_io_out_0_bits_25),
    .io_out_0_bits_26(aluOutputDemux_x6_demux_io_out_0_bits_26),
    .io_out_0_bits_27(aluOutputDemux_x6_demux_io_out_0_bits_27),
    .io_out_0_bits_28(aluOutputDemux_x6_demux_io_out_0_bits_28),
    .io_out_0_bits_29(aluOutputDemux_x6_demux_io_out_0_bits_29),
    .io_out_0_bits_30(aluOutputDemux_x6_demux_io_out_0_bits_30),
    .io_out_0_bits_31(aluOutputDemux_x6_demux_io_out_0_bits_31),
    .io_out_1_ready(aluOutputDemux_x6_demux_io_out_1_ready),
    .io_out_1_valid(aluOutputDemux_x6_demux_io_out_1_valid),
    .io_out_1_bits_0(aluOutputDemux_x6_demux_io_out_1_bits_0),
    .io_out_1_bits_1(aluOutputDemux_x6_demux_io_out_1_bits_1),
    .io_out_1_bits_2(aluOutputDemux_x6_demux_io_out_1_bits_2),
    .io_out_1_bits_3(aluOutputDemux_x6_demux_io_out_1_bits_3),
    .io_out_1_bits_4(aluOutputDemux_x6_demux_io_out_1_bits_4),
    .io_out_1_bits_5(aluOutputDemux_x6_demux_io_out_1_bits_5),
    .io_out_1_bits_6(aluOutputDemux_x6_demux_io_out_1_bits_6),
    .io_out_1_bits_7(aluOutputDemux_x6_demux_io_out_1_bits_7),
    .io_out_1_bits_8(aluOutputDemux_x6_demux_io_out_1_bits_8),
    .io_out_1_bits_9(aluOutputDemux_x6_demux_io_out_1_bits_9),
    .io_out_1_bits_10(aluOutputDemux_x6_demux_io_out_1_bits_10),
    .io_out_1_bits_11(aluOutputDemux_x6_demux_io_out_1_bits_11),
    .io_out_1_bits_12(aluOutputDemux_x6_demux_io_out_1_bits_12),
    .io_out_1_bits_13(aluOutputDemux_x6_demux_io_out_1_bits_13),
    .io_out_1_bits_14(aluOutputDemux_x6_demux_io_out_1_bits_14),
    .io_out_1_bits_15(aluOutputDemux_x6_demux_io_out_1_bits_15),
    .io_out_1_bits_16(aluOutputDemux_x6_demux_io_out_1_bits_16),
    .io_out_1_bits_17(aluOutputDemux_x6_demux_io_out_1_bits_17),
    .io_out_1_bits_18(aluOutputDemux_x6_demux_io_out_1_bits_18),
    .io_out_1_bits_19(aluOutputDemux_x6_demux_io_out_1_bits_19),
    .io_out_1_bits_20(aluOutputDemux_x6_demux_io_out_1_bits_20),
    .io_out_1_bits_21(aluOutputDemux_x6_demux_io_out_1_bits_21),
    .io_out_1_bits_22(aluOutputDemux_x6_demux_io_out_1_bits_22),
    .io_out_1_bits_23(aluOutputDemux_x6_demux_io_out_1_bits_23),
    .io_out_1_bits_24(aluOutputDemux_x6_demux_io_out_1_bits_24),
    .io_out_1_bits_25(aluOutputDemux_x6_demux_io_out_1_bits_25),
    .io_out_1_bits_26(aluOutputDemux_x6_demux_io_out_1_bits_26),
    .io_out_1_bits_27(aluOutputDemux_x6_demux_io_out_1_bits_27),
    .io_out_1_bits_28(aluOutputDemux_x6_demux_io_out_1_bits_28),
    .io_out_1_bits_29(aluOutputDemux_x6_demux_io_out_1_bits_29),
    .io_out_1_bits_30(aluOutputDemux_x6_demux_io_out_1_bits_30),
    .io_out_1_bits_31(aluOutputDemux_x6_demux_io_out_1_bits_31)
  );
  Queue_15 aluOutputDemux ( // @[Mem.scala 22:19]
    .clock(aluOutputDemux_clock),
    .reset(aluOutputDemux_reset),
    .io_enq_ready(aluOutputDemux_io_enq_ready),
    .io_enq_valid(aluOutputDemux_io_enq_valid),
    .io_enq_bits(aluOutputDemux_io_enq_bits),
    .io_deq_ready(aluOutputDemux_io_deq_ready),
    .io_deq_valid(aluOutputDemux_io_deq_valid),
    .io_deq_bits(aluOutputDemux_io_deq_bits)
  );
  Mux accInputMux_x15_mux ( // @[Mux.scala 71:21]
    .io_in_0_ready(accInputMux_x15_mux_io_in_0_ready),
    .io_in_0_valid(accInputMux_x15_mux_io_in_0_valid),
    .io_in_0_bits_0(accInputMux_x15_mux_io_in_0_bits_0),
    .io_in_0_bits_1(accInputMux_x15_mux_io_in_0_bits_1),
    .io_in_0_bits_2(accInputMux_x15_mux_io_in_0_bits_2),
    .io_in_0_bits_3(accInputMux_x15_mux_io_in_0_bits_3),
    .io_in_0_bits_4(accInputMux_x15_mux_io_in_0_bits_4),
    .io_in_0_bits_5(accInputMux_x15_mux_io_in_0_bits_5),
    .io_in_0_bits_6(accInputMux_x15_mux_io_in_0_bits_6),
    .io_in_0_bits_7(accInputMux_x15_mux_io_in_0_bits_7),
    .io_in_0_bits_8(accInputMux_x15_mux_io_in_0_bits_8),
    .io_in_0_bits_9(accInputMux_x15_mux_io_in_0_bits_9),
    .io_in_0_bits_10(accInputMux_x15_mux_io_in_0_bits_10),
    .io_in_0_bits_11(accInputMux_x15_mux_io_in_0_bits_11),
    .io_in_0_bits_12(accInputMux_x15_mux_io_in_0_bits_12),
    .io_in_0_bits_13(accInputMux_x15_mux_io_in_0_bits_13),
    .io_in_0_bits_14(accInputMux_x15_mux_io_in_0_bits_14),
    .io_in_0_bits_15(accInputMux_x15_mux_io_in_0_bits_15),
    .io_in_0_bits_16(accInputMux_x15_mux_io_in_0_bits_16),
    .io_in_0_bits_17(accInputMux_x15_mux_io_in_0_bits_17),
    .io_in_0_bits_18(accInputMux_x15_mux_io_in_0_bits_18),
    .io_in_0_bits_19(accInputMux_x15_mux_io_in_0_bits_19),
    .io_in_0_bits_20(accInputMux_x15_mux_io_in_0_bits_20),
    .io_in_0_bits_21(accInputMux_x15_mux_io_in_0_bits_21),
    .io_in_0_bits_22(accInputMux_x15_mux_io_in_0_bits_22),
    .io_in_0_bits_23(accInputMux_x15_mux_io_in_0_bits_23),
    .io_in_0_bits_24(accInputMux_x15_mux_io_in_0_bits_24),
    .io_in_0_bits_25(accInputMux_x15_mux_io_in_0_bits_25),
    .io_in_0_bits_26(accInputMux_x15_mux_io_in_0_bits_26),
    .io_in_0_bits_27(accInputMux_x15_mux_io_in_0_bits_27),
    .io_in_0_bits_28(accInputMux_x15_mux_io_in_0_bits_28),
    .io_in_0_bits_29(accInputMux_x15_mux_io_in_0_bits_29),
    .io_in_0_bits_30(accInputMux_x15_mux_io_in_0_bits_30),
    .io_in_0_bits_31(accInputMux_x15_mux_io_in_0_bits_31),
    .io_in_1_ready(accInputMux_x15_mux_io_in_1_ready),
    .io_in_1_valid(accInputMux_x15_mux_io_in_1_valid),
    .io_in_1_bits_0(accInputMux_x15_mux_io_in_1_bits_0),
    .io_in_1_bits_1(accInputMux_x15_mux_io_in_1_bits_1),
    .io_in_1_bits_2(accInputMux_x15_mux_io_in_1_bits_2),
    .io_in_1_bits_3(accInputMux_x15_mux_io_in_1_bits_3),
    .io_in_1_bits_4(accInputMux_x15_mux_io_in_1_bits_4),
    .io_in_1_bits_5(accInputMux_x15_mux_io_in_1_bits_5),
    .io_in_1_bits_6(accInputMux_x15_mux_io_in_1_bits_6),
    .io_in_1_bits_7(accInputMux_x15_mux_io_in_1_bits_7),
    .io_in_1_bits_8(accInputMux_x15_mux_io_in_1_bits_8),
    .io_in_1_bits_9(accInputMux_x15_mux_io_in_1_bits_9),
    .io_in_1_bits_10(accInputMux_x15_mux_io_in_1_bits_10),
    .io_in_1_bits_11(accInputMux_x15_mux_io_in_1_bits_11),
    .io_in_1_bits_12(accInputMux_x15_mux_io_in_1_bits_12),
    .io_in_1_bits_13(accInputMux_x15_mux_io_in_1_bits_13),
    .io_in_1_bits_14(accInputMux_x15_mux_io_in_1_bits_14),
    .io_in_1_bits_15(accInputMux_x15_mux_io_in_1_bits_15),
    .io_in_1_bits_16(accInputMux_x15_mux_io_in_1_bits_16),
    .io_in_1_bits_17(accInputMux_x15_mux_io_in_1_bits_17),
    .io_in_1_bits_18(accInputMux_x15_mux_io_in_1_bits_18),
    .io_in_1_bits_19(accInputMux_x15_mux_io_in_1_bits_19),
    .io_in_1_bits_20(accInputMux_x15_mux_io_in_1_bits_20),
    .io_in_1_bits_21(accInputMux_x15_mux_io_in_1_bits_21),
    .io_in_1_bits_22(accInputMux_x15_mux_io_in_1_bits_22),
    .io_in_1_bits_23(accInputMux_x15_mux_io_in_1_bits_23),
    .io_in_1_bits_24(accInputMux_x15_mux_io_in_1_bits_24),
    .io_in_1_bits_25(accInputMux_x15_mux_io_in_1_bits_25),
    .io_in_1_bits_26(accInputMux_x15_mux_io_in_1_bits_26),
    .io_in_1_bits_27(accInputMux_x15_mux_io_in_1_bits_27),
    .io_in_1_bits_28(accInputMux_x15_mux_io_in_1_bits_28),
    .io_in_1_bits_29(accInputMux_x15_mux_io_in_1_bits_29),
    .io_in_1_bits_30(accInputMux_x15_mux_io_in_1_bits_30),
    .io_in_1_bits_31(accInputMux_x15_mux_io_in_1_bits_31),
    .io_sel_ready(accInputMux_x15_mux_io_sel_ready),
    .io_sel_valid(accInputMux_x15_mux_io_sel_valid),
    .io_sel_bits(accInputMux_x15_mux_io_sel_bits),
    .io_out_ready(accInputMux_x15_mux_io_out_ready),
    .io_out_valid(accInputMux_x15_mux_io_out_valid),
    .io_out_bits_0(accInputMux_x15_mux_io_out_bits_0),
    .io_out_bits_1(accInputMux_x15_mux_io_out_bits_1),
    .io_out_bits_2(accInputMux_x15_mux_io_out_bits_2),
    .io_out_bits_3(accInputMux_x15_mux_io_out_bits_3),
    .io_out_bits_4(accInputMux_x15_mux_io_out_bits_4),
    .io_out_bits_5(accInputMux_x15_mux_io_out_bits_5),
    .io_out_bits_6(accInputMux_x15_mux_io_out_bits_6),
    .io_out_bits_7(accInputMux_x15_mux_io_out_bits_7),
    .io_out_bits_8(accInputMux_x15_mux_io_out_bits_8),
    .io_out_bits_9(accInputMux_x15_mux_io_out_bits_9),
    .io_out_bits_10(accInputMux_x15_mux_io_out_bits_10),
    .io_out_bits_11(accInputMux_x15_mux_io_out_bits_11),
    .io_out_bits_12(accInputMux_x15_mux_io_out_bits_12),
    .io_out_bits_13(accInputMux_x15_mux_io_out_bits_13),
    .io_out_bits_14(accInputMux_x15_mux_io_out_bits_14),
    .io_out_bits_15(accInputMux_x15_mux_io_out_bits_15),
    .io_out_bits_16(accInputMux_x15_mux_io_out_bits_16),
    .io_out_bits_17(accInputMux_x15_mux_io_out_bits_17),
    .io_out_bits_18(accInputMux_x15_mux_io_out_bits_18),
    .io_out_bits_19(accInputMux_x15_mux_io_out_bits_19),
    .io_out_bits_20(accInputMux_x15_mux_io_out_bits_20),
    .io_out_bits_21(accInputMux_x15_mux_io_out_bits_21),
    .io_out_bits_22(accInputMux_x15_mux_io_out_bits_22),
    .io_out_bits_23(accInputMux_x15_mux_io_out_bits_23),
    .io_out_bits_24(accInputMux_x15_mux_io_out_bits_24),
    .io_out_bits_25(accInputMux_x15_mux_io_out_bits_25),
    .io_out_bits_26(accInputMux_x15_mux_io_out_bits_26),
    .io_out_bits_27(accInputMux_x15_mux_io_out_bits_27),
    .io_out_bits_28(accInputMux_x15_mux_io_out_bits_28),
    .io_out_bits_29(accInputMux_x15_mux_io_out_bits_29),
    .io_out_bits_30(accInputMux_x15_mux_io_out_bits_30),
    .io_out_bits_31(accInputMux_x15_mux_io_out_bits_31)
  );
  Queue_15 accInputMux ( // @[Mem.scala 22:19]
    .clock(accInputMux_clock),
    .reset(accInputMux_reset),
    .io_enq_ready(accInputMux_io_enq_ready),
    .io_enq_valid(accInputMux_io_enq_valid),
    .io_enq_bits(accInputMux_io_enq_bits),
    .io_deq_ready(accInputMux_io_deq_ready),
    .io_deq_valid(accInputMux_io_deq_valid),
    .io_deq_bits(accInputMux_io_deq_bits)
  );
  Demux accOutputDemux_x24_demux ( // @[Demux.scala 46:23]
    .io_in_ready(accOutputDemux_x24_demux_io_in_ready),
    .io_in_valid(accOutputDemux_x24_demux_io_in_valid),
    .io_in_bits_0(accOutputDemux_x24_demux_io_in_bits_0),
    .io_in_bits_1(accOutputDemux_x24_demux_io_in_bits_1),
    .io_in_bits_2(accOutputDemux_x24_demux_io_in_bits_2),
    .io_in_bits_3(accOutputDemux_x24_demux_io_in_bits_3),
    .io_in_bits_4(accOutputDemux_x24_demux_io_in_bits_4),
    .io_in_bits_5(accOutputDemux_x24_demux_io_in_bits_5),
    .io_in_bits_6(accOutputDemux_x24_demux_io_in_bits_6),
    .io_in_bits_7(accOutputDemux_x24_demux_io_in_bits_7),
    .io_in_bits_8(accOutputDemux_x24_demux_io_in_bits_8),
    .io_in_bits_9(accOutputDemux_x24_demux_io_in_bits_9),
    .io_in_bits_10(accOutputDemux_x24_demux_io_in_bits_10),
    .io_in_bits_11(accOutputDemux_x24_demux_io_in_bits_11),
    .io_in_bits_12(accOutputDemux_x24_demux_io_in_bits_12),
    .io_in_bits_13(accOutputDemux_x24_demux_io_in_bits_13),
    .io_in_bits_14(accOutputDemux_x24_demux_io_in_bits_14),
    .io_in_bits_15(accOutputDemux_x24_demux_io_in_bits_15),
    .io_in_bits_16(accOutputDemux_x24_demux_io_in_bits_16),
    .io_in_bits_17(accOutputDemux_x24_demux_io_in_bits_17),
    .io_in_bits_18(accOutputDemux_x24_demux_io_in_bits_18),
    .io_in_bits_19(accOutputDemux_x24_demux_io_in_bits_19),
    .io_in_bits_20(accOutputDemux_x24_demux_io_in_bits_20),
    .io_in_bits_21(accOutputDemux_x24_demux_io_in_bits_21),
    .io_in_bits_22(accOutputDemux_x24_demux_io_in_bits_22),
    .io_in_bits_23(accOutputDemux_x24_demux_io_in_bits_23),
    .io_in_bits_24(accOutputDemux_x24_demux_io_in_bits_24),
    .io_in_bits_25(accOutputDemux_x24_demux_io_in_bits_25),
    .io_in_bits_26(accOutputDemux_x24_demux_io_in_bits_26),
    .io_in_bits_27(accOutputDemux_x24_demux_io_in_bits_27),
    .io_in_bits_28(accOutputDemux_x24_demux_io_in_bits_28),
    .io_in_bits_29(accOutputDemux_x24_demux_io_in_bits_29),
    .io_in_bits_30(accOutputDemux_x24_demux_io_in_bits_30),
    .io_in_bits_31(accOutputDemux_x24_demux_io_in_bits_31),
    .io_sel_ready(accOutputDemux_x24_demux_io_sel_ready),
    .io_sel_valid(accOutputDemux_x24_demux_io_sel_valid),
    .io_sel_bits(accOutputDemux_x24_demux_io_sel_bits),
    .io_out_0_ready(accOutputDemux_x24_demux_io_out_0_ready),
    .io_out_0_valid(accOutputDemux_x24_demux_io_out_0_valid),
    .io_out_0_bits_0(accOutputDemux_x24_demux_io_out_0_bits_0),
    .io_out_0_bits_1(accOutputDemux_x24_demux_io_out_0_bits_1),
    .io_out_0_bits_2(accOutputDemux_x24_demux_io_out_0_bits_2),
    .io_out_0_bits_3(accOutputDemux_x24_demux_io_out_0_bits_3),
    .io_out_0_bits_4(accOutputDemux_x24_demux_io_out_0_bits_4),
    .io_out_0_bits_5(accOutputDemux_x24_demux_io_out_0_bits_5),
    .io_out_0_bits_6(accOutputDemux_x24_demux_io_out_0_bits_6),
    .io_out_0_bits_7(accOutputDemux_x24_demux_io_out_0_bits_7),
    .io_out_0_bits_8(accOutputDemux_x24_demux_io_out_0_bits_8),
    .io_out_0_bits_9(accOutputDemux_x24_demux_io_out_0_bits_9),
    .io_out_0_bits_10(accOutputDemux_x24_demux_io_out_0_bits_10),
    .io_out_0_bits_11(accOutputDemux_x24_demux_io_out_0_bits_11),
    .io_out_0_bits_12(accOutputDemux_x24_demux_io_out_0_bits_12),
    .io_out_0_bits_13(accOutputDemux_x24_demux_io_out_0_bits_13),
    .io_out_0_bits_14(accOutputDemux_x24_demux_io_out_0_bits_14),
    .io_out_0_bits_15(accOutputDemux_x24_demux_io_out_0_bits_15),
    .io_out_0_bits_16(accOutputDemux_x24_demux_io_out_0_bits_16),
    .io_out_0_bits_17(accOutputDemux_x24_demux_io_out_0_bits_17),
    .io_out_0_bits_18(accOutputDemux_x24_demux_io_out_0_bits_18),
    .io_out_0_bits_19(accOutputDemux_x24_demux_io_out_0_bits_19),
    .io_out_0_bits_20(accOutputDemux_x24_demux_io_out_0_bits_20),
    .io_out_0_bits_21(accOutputDemux_x24_demux_io_out_0_bits_21),
    .io_out_0_bits_22(accOutputDemux_x24_demux_io_out_0_bits_22),
    .io_out_0_bits_23(accOutputDemux_x24_demux_io_out_0_bits_23),
    .io_out_0_bits_24(accOutputDemux_x24_demux_io_out_0_bits_24),
    .io_out_0_bits_25(accOutputDemux_x24_demux_io_out_0_bits_25),
    .io_out_0_bits_26(accOutputDemux_x24_demux_io_out_0_bits_26),
    .io_out_0_bits_27(accOutputDemux_x24_demux_io_out_0_bits_27),
    .io_out_0_bits_28(accOutputDemux_x24_demux_io_out_0_bits_28),
    .io_out_0_bits_29(accOutputDemux_x24_demux_io_out_0_bits_29),
    .io_out_0_bits_30(accOutputDemux_x24_demux_io_out_0_bits_30),
    .io_out_0_bits_31(accOutputDemux_x24_demux_io_out_0_bits_31),
    .io_out_1_ready(accOutputDemux_x24_demux_io_out_1_ready),
    .io_out_1_valid(accOutputDemux_x24_demux_io_out_1_valid),
    .io_out_1_bits_0(accOutputDemux_x24_demux_io_out_1_bits_0),
    .io_out_1_bits_1(accOutputDemux_x24_demux_io_out_1_bits_1),
    .io_out_1_bits_2(accOutputDemux_x24_demux_io_out_1_bits_2),
    .io_out_1_bits_3(accOutputDemux_x24_demux_io_out_1_bits_3),
    .io_out_1_bits_4(accOutputDemux_x24_demux_io_out_1_bits_4),
    .io_out_1_bits_5(accOutputDemux_x24_demux_io_out_1_bits_5),
    .io_out_1_bits_6(accOutputDemux_x24_demux_io_out_1_bits_6),
    .io_out_1_bits_7(accOutputDemux_x24_demux_io_out_1_bits_7),
    .io_out_1_bits_8(accOutputDemux_x24_demux_io_out_1_bits_8),
    .io_out_1_bits_9(accOutputDemux_x24_demux_io_out_1_bits_9),
    .io_out_1_bits_10(accOutputDemux_x24_demux_io_out_1_bits_10),
    .io_out_1_bits_11(accOutputDemux_x24_demux_io_out_1_bits_11),
    .io_out_1_bits_12(accOutputDemux_x24_demux_io_out_1_bits_12),
    .io_out_1_bits_13(accOutputDemux_x24_demux_io_out_1_bits_13),
    .io_out_1_bits_14(accOutputDemux_x24_demux_io_out_1_bits_14),
    .io_out_1_bits_15(accOutputDemux_x24_demux_io_out_1_bits_15),
    .io_out_1_bits_16(accOutputDemux_x24_demux_io_out_1_bits_16),
    .io_out_1_bits_17(accOutputDemux_x24_demux_io_out_1_bits_17),
    .io_out_1_bits_18(accOutputDemux_x24_demux_io_out_1_bits_18),
    .io_out_1_bits_19(accOutputDemux_x24_demux_io_out_1_bits_19),
    .io_out_1_bits_20(accOutputDemux_x24_demux_io_out_1_bits_20),
    .io_out_1_bits_21(accOutputDemux_x24_demux_io_out_1_bits_21),
    .io_out_1_bits_22(accOutputDemux_x24_demux_io_out_1_bits_22),
    .io_out_1_bits_23(accOutputDemux_x24_demux_io_out_1_bits_23),
    .io_out_1_bits_24(accOutputDemux_x24_demux_io_out_1_bits_24),
    .io_out_1_bits_25(accOutputDemux_x24_demux_io_out_1_bits_25),
    .io_out_1_bits_26(accOutputDemux_x24_demux_io_out_1_bits_26),
    .io_out_1_bits_27(accOutputDemux_x24_demux_io_out_1_bits_27),
    .io_out_1_bits_28(accOutputDemux_x24_demux_io_out_1_bits_28),
    .io_out_1_bits_29(accOutputDemux_x24_demux_io_out_1_bits_29),
    .io_out_1_bits_30(accOutputDemux_x24_demux_io_out_1_bits_30),
    .io_out_1_bits_31(accOutputDemux_x24_demux_io_out_1_bits_31)
  );
  Queue_15 accOutputDemux ( // @[Mem.scala 22:19]
    .clock(accOutputDemux_clock),
    .reset(accOutputDemux_reset),
    .io_enq_ready(accOutputDemux_io_enq_ready),
    .io_enq_valid(accOutputDemux_io_enq_valid),
    .io_enq_bits(accOutputDemux_io_enq_bits),
    .io_deq_ready(accOutputDemux_io_deq_ready),
    .io_deq_valid(accOutputDemux_io_deq_valid),
    .io_deq_bits(accOutputDemux_io_deq_bits)
  );
  MultiEnqueue_1 accWriteEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(accWriteEnqueuer_clock),
    .reset(accWriteEnqueuer_reset),
    .io_in_ready(accWriteEnqueuer_io_in_ready),
    .io_in_valid(accWriteEnqueuer_io_in_valid),
    .io_out_0_ready(accWriteEnqueuer_io_out_0_ready),
    .io_out_0_valid(accWriteEnqueuer_io_out_0_valid),
    .io_out_1_ready(accWriteEnqueuer_io_out_1_ready),
    .io_out_1_valid(accWriteEnqueuer_io_out_1_valid)
  );
  MultiEnqueue_1 accReadEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(accReadEnqueuer_clock),
    .reset(accReadEnqueuer_reset),
    .io_in_ready(accReadEnqueuer_io_in_ready),
    .io_in_valid(accReadEnqueuer_io_in_valid),
    .io_out_0_ready(accReadEnqueuer_io_out_0_ready),
    .io_out_0_valid(accReadEnqueuer_io_out_0_valid),
    .io_out_1_ready(accReadEnqueuer_io_out_1_ready),
    .io_out_1_valid(accReadEnqueuer_io_out_1_valid)
  );
  MultiEnqueue_2 simdRWWriteEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(simdRWWriteEnqueuer_clock),
    .reset(simdRWWriteEnqueuer_reset),
    .io_in_ready(simdRWWriteEnqueuer_io_in_ready),
    .io_in_valid(simdRWWriteEnqueuer_io_in_valid),
    .io_out_0_ready(simdRWWriteEnqueuer_io_out_0_ready),
    .io_out_0_valid(simdRWWriteEnqueuer_io_out_0_valid),
    .io_out_1_ready(simdRWWriteEnqueuer_io_out_1_ready),
    .io_out_1_valid(simdRWWriteEnqueuer_io_out_1_valid),
    .io_out_2_ready(simdRWWriteEnqueuer_io_out_2_ready),
    .io_out_2_valid(simdRWWriteEnqueuer_io_out_2_valid)
  );
  MultiEnqueue_2 simdRWReadEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(simdRWReadEnqueuer_clock),
    .reset(simdRWReadEnqueuer_reset),
    .io_in_ready(simdRWReadEnqueuer_io_in_ready),
    .io_in_valid(simdRWReadEnqueuer_io_in_valid),
    .io_out_0_ready(simdRWReadEnqueuer_io_out_0_ready),
    .io_out_0_valid(simdRWReadEnqueuer_io_out_0_valid),
    .io_out_1_ready(simdRWReadEnqueuer_io_out_1_ready),
    .io_out_1_valid(simdRWReadEnqueuer_io_out_1_valid),
    .io_out_2_ready(simdRWReadEnqueuer_io_out_2_ready),
    .io_out_2_valid(simdRWReadEnqueuer_io_out_2_valid)
  );
  MultiEnqueue_3 simdWriteEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(simdWriteEnqueuer_clock),
    .reset(simdWriteEnqueuer_reset),
    .io_in_ready(simdWriteEnqueuer_io_in_ready),
    .io_in_valid(simdWriteEnqueuer_io_in_valid),
    .io_out_0_ready(simdWriteEnqueuer_io_out_0_ready),
    .io_out_0_valid(simdWriteEnqueuer_io_out_0_valid),
    .io_out_1_ready(simdWriteEnqueuer_io_out_1_ready),
    .io_out_1_valid(simdWriteEnqueuer_io_out_1_valid),
    .io_out_2_ready(simdWriteEnqueuer_io_out_2_ready),
    .io_out_2_valid(simdWriteEnqueuer_io_out_2_valid),
    .io_out_3_ready(simdWriteEnqueuer_io_out_3_ready),
    .io_out_3_valid(simdWriteEnqueuer_io_out_3_valid)
  );
  MultiEnqueue_3 simdReadEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(simdReadEnqueuer_clock),
    .reset(simdReadEnqueuer_reset),
    .io_in_ready(simdReadEnqueuer_io_in_ready),
    .io_in_valid(simdReadEnqueuer_io_in_valid),
    .io_out_0_ready(simdReadEnqueuer_io_out_0_ready),
    .io_out_0_valid(simdReadEnqueuer_io_out_0_valid),
    .io_out_1_ready(simdReadEnqueuer_io_out_1_ready),
    .io_out_1_valid(simdReadEnqueuer_io_out_1_valid),
    .io_out_2_ready(simdReadEnqueuer_io_out_2_ready),
    .io_out_2_valid(simdReadEnqueuer_io_out_2_valid),
    .io_out_3_ready(simdReadEnqueuer_io_out_3_ready),
    .io_out_3_valid(simdReadEnqueuer_io_out_3_valid)
  );
  MultiEnqueue_1 simdEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(simdEnqueuer_clock),
    .reset(simdEnqueuer_reset),
    .io_in_ready(simdEnqueuer_io_in_ready),
    .io_in_valid(simdEnqueuer_io_in_valid),
    .io_out_0_ready(simdEnqueuer_io_out_0_ready),
    .io_out_0_valid(simdEnqueuer_io_out_0_valid),
    .io_out_1_ready(simdEnqueuer_io_out_1_ready),
    .io_out_1_valid(simdEnqueuer_io_out_1_valid)
  );
  assign io_input_ready = accInputMux_x15_mux_io_in_0_ready; // @[Mux.scala 79:18]
  assign io_output_valid = accOutputDemux_x24_demux_io_out_0_valid; // @[Demux.scala 55:10]
  assign io_output_bits_0 = accOutputDemux_x24_demux_io_out_0_bits_0; // @[Demux.scala 55:10]
  assign io_output_bits_1 = accOutputDemux_x24_demux_io_out_0_bits_1; // @[Demux.scala 55:10]
  assign io_output_bits_2 = accOutputDemux_x24_demux_io_out_0_bits_2; // @[Demux.scala 55:10]
  assign io_output_bits_3 = accOutputDemux_x24_demux_io_out_0_bits_3; // @[Demux.scala 55:10]
  assign io_output_bits_4 = accOutputDemux_x24_demux_io_out_0_bits_4; // @[Demux.scala 55:10]
  assign io_output_bits_5 = accOutputDemux_x24_demux_io_out_0_bits_5; // @[Demux.scala 55:10]
  assign io_output_bits_6 = accOutputDemux_x24_demux_io_out_0_bits_6; // @[Demux.scala 55:10]
  assign io_output_bits_7 = accOutputDemux_x24_demux_io_out_0_bits_7; // @[Demux.scala 55:10]
  assign io_output_bits_8 = accOutputDemux_x24_demux_io_out_0_bits_8; // @[Demux.scala 55:10]
  assign io_output_bits_9 = accOutputDemux_x24_demux_io_out_0_bits_9; // @[Demux.scala 55:10]
  assign io_output_bits_10 = accOutputDemux_x24_demux_io_out_0_bits_10; // @[Demux.scala 55:10]
  assign io_output_bits_11 = accOutputDemux_x24_demux_io_out_0_bits_11; // @[Demux.scala 55:10]
  assign io_output_bits_12 = accOutputDemux_x24_demux_io_out_0_bits_12; // @[Demux.scala 55:10]
  assign io_output_bits_13 = accOutputDemux_x24_demux_io_out_0_bits_13; // @[Demux.scala 55:10]
  assign io_output_bits_14 = accOutputDemux_x24_demux_io_out_0_bits_14; // @[Demux.scala 55:10]
  assign io_output_bits_15 = accOutputDemux_x24_demux_io_out_0_bits_15; // @[Demux.scala 55:10]
  assign io_output_bits_16 = accOutputDemux_x24_demux_io_out_0_bits_16; // @[Demux.scala 55:10]
  assign io_output_bits_17 = accOutputDemux_x24_demux_io_out_0_bits_17; // @[Demux.scala 55:10]
  assign io_output_bits_18 = accOutputDemux_x24_demux_io_out_0_bits_18; // @[Demux.scala 55:10]
  assign io_output_bits_19 = accOutputDemux_x24_demux_io_out_0_bits_19; // @[Demux.scala 55:10]
  assign io_output_bits_20 = accOutputDemux_x24_demux_io_out_0_bits_20; // @[Demux.scala 55:10]
  assign io_output_bits_21 = accOutputDemux_x24_demux_io_out_0_bits_21; // @[Demux.scala 55:10]
  assign io_output_bits_22 = accOutputDemux_x24_demux_io_out_0_bits_22; // @[Demux.scala 55:10]
  assign io_output_bits_23 = accOutputDemux_x24_demux_io_out_0_bits_23; // @[Demux.scala 55:10]
  assign io_output_bits_24 = accOutputDemux_x24_demux_io_out_0_bits_24; // @[Demux.scala 55:10]
  assign io_output_bits_25 = accOutputDemux_x24_demux_io_out_0_bits_25; // @[Demux.scala 55:10]
  assign io_output_bits_26 = accOutputDemux_x24_demux_io_out_0_bits_26; // @[Demux.scala 55:10]
  assign io_output_bits_27 = accOutputDemux_x24_demux_io_out_0_bits_27; // @[Demux.scala 55:10]
  assign io_output_bits_28 = accOutputDemux_x24_demux_io_out_0_bits_28; // @[Demux.scala 55:10]
  assign io_output_bits_29 = accOutputDemux_x24_demux_io_out_0_bits_29; // @[Demux.scala 55:10]
  assign io_output_bits_30 = accOutputDemux_x24_demux_io_out_0_bits_30; // @[Demux.scala 55:10]
  assign io_output_bits_31 = accOutputDemux_x24_demux_io_out_0_bits_31; // @[Demux.scala 55:10]
  assign io_control_ready = isNoOp ? dataPathReady : dataPathReady_1; // @[AccumulatorWithALUArray.scala 133:16 182:19 257:19]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_io_input_valid = accInputMux_x15_mux_io_out_valid; // @[Mux.scala 81:9]
  assign acc_io_input_bits_0 = accInputMux_x15_mux_io_out_bits_0; // @[Mux.scala 81:9]
  assign acc_io_input_bits_1 = accInputMux_x15_mux_io_out_bits_1; // @[Mux.scala 81:9]
  assign acc_io_input_bits_2 = accInputMux_x15_mux_io_out_bits_2; // @[Mux.scala 81:9]
  assign acc_io_input_bits_3 = accInputMux_x15_mux_io_out_bits_3; // @[Mux.scala 81:9]
  assign acc_io_input_bits_4 = accInputMux_x15_mux_io_out_bits_4; // @[Mux.scala 81:9]
  assign acc_io_input_bits_5 = accInputMux_x15_mux_io_out_bits_5; // @[Mux.scala 81:9]
  assign acc_io_input_bits_6 = accInputMux_x15_mux_io_out_bits_6; // @[Mux.scala 81:9]
  assign acc_io_input_bits_7 = accInputMux_x15_mux_io_out_bits_7; // @[Mux.scala 81:9]
  assign acc_io_input_bits_8 = accInputMux_x15_mux_io_out_bits_8; // @[Mux.scala 81:9]
  assign acc_io_input_bits_9 = accInputMux_x15_mux_io_out_bits_9; // @[Mux.scala 81:9]
  assign acc_io_input_bits_10 = accInputMux_x15_mux_io_out_bits_10; // @[Mux.scala 81:9]
  assign acc_io_input_bits_11 = accInputMux_x15_mux_io_out_bits_11; // @[Mux.scala 81:9]
  assign acc_io_input_bits_12 = accInputMux_x15_mux_io_out_bits_12; // @[Mux.scala 81:9]
  assign acc_io_input_bits_13 = accInputMux_x15_mux_io_out_bits_13; // @[Mux.scala 81:9]
  assign acc_io_input_bits_14 = accInputMux_x15_mux_io_out_bits_14; // @[Mux.scala 81:9]
  assign acc_io_input_bits_15 = accInputMux_x15_mux_io_out_bits_15; // @[Mux.scala 81:9]
  assign acc_io_input_bits_16 = accInputMux_x15_mux_io_out_bits_16; // @[Mux.scala 81:9]
  assign acc_io_input_bits_17 = accInputMux_x15_mux_io_out_bits_17; // @[Mux.scala 81:9]
  assign acc_io_input_bits_18 = accInputMux_x15_mux_io_out_bits_18; // @[Mux.scala 81:9]
  assign acc_io_input_bits_19 = accInputMux_x15_mux_io_out_bits_19; // @[Mux.scala 81:9]
  assign acc_io_input_bits_20 = accInputMux_x15_mux_io_out_bits_20; // @[Mux.scala 81:9]
  assign acc_io_input_bits_21 = accInputMux_x15_mux_io_out_bits_21; // @[Mux.scala 81:9]
  assign acc_io_input_bits_22 = accInputMux_x15_mux_io_out_bits_22; // @[Mux.scala 81:9]
  assign acc_io_input_bits_23 = accInputMux_x15_mux_io_out_bits_23; // @[Mux.scala 81:9]
  assign acc_io_input_bits_24 = accInputMux_x15_mux_io_out_bits_24; // @[Mux.scala 81:9]
  assign acc_io_input_bits_25 = accInputMux_x15_mux_io_out_bits_25; // @[Mux.scala 81:9]
  assign acc_io_input_bits_26 = accInputMux_x15_mux_io_out_bits_26; // @[Mux.scala 81:9]
  assign acc_io_input_bits_27 = accInputMux_x15_mux_io_out_bits_27; // @[Mux.scala 81:9]
  assign acc_io_input_bits_28 = accInputMux_x15_mux_io_out_bits_28; // @[Mux.scala 81:9]
  assign acc_io_input_bits_29 = accInputMux_x15_mux_io_out_bits_29; // @[Mux.scala 81:9]
  assign acc_io_input_bits_30 = accInputMux_x15_mux_io_out_bits_30; // @[Mux.scala 81:9]
  assign acc_io_input_bits_31 = accInputMux_x15_mux_io_out_bits_31; // @[Mux.scala 81:9]
  assign acc_io_output_ready = accOutputDemux_x24_demux_io_in_ready; // @[Demux.scala 54:17]
  assign acc_io_control_valid = isNoOp ? _GEN_45 : _GEN_151; // @[AccumulatorWithALUArray.scala 133:16]
  assign acc_io_control_bits_address = isNoOp ? _GEN_46 : _GEN_152; // @[AccumulatorWithALUArray.scala 133:16]
  assign acc_io_control_bits_accumulate = isNoOp ? _GEN_47 : _GEN_47; // @[AccumulatorWithALUArray.scala 133:16]
  assign acc_io_control_bits_write = isNoOp ? _GEN_48 : _GEN_48; // @[AccumulatorWithALUArray.scala 133:16]
  assign acc_io_tracepoint = io_tracepoint; // @[AccumulatorWithALUArray.scala 68:21]
  assign acc_io_programCounter = io_programCounter; // @[AccumulatorWithALUArray.scala 69:25]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_input_valid = accOutputDemux_x24_demux_io_out_1_valid; // @[Demux.scala 56:10]
  assign alu_io_input_bits_0 = accOutputDemux_x24_demux_io_out_1_bits_0; // @[Demux.scala 56:10]
  assign alu_io_input_bits_1 = accOutputDemux_x24_demux_io_out_1_bits_1; // @[Demux.scala 56:10]
  assign alu_io_input_bits_2 = accOutputDemux_x24_demux_io_out_1_bits_2; // @[Demux.scala 56:10]
  assign alu_io_input_bits_3 = accOutputDemux_x24_demux_io_out_1_bits_3; // @[Demux.scala 56:10]
  assign alu_io_input_bits_4 = accOutputDemux_x24_demux_io_out_1_bits_4; // @[Demux.scala 56:10]
  assign alu_io_input_bits_5 = accOutputDemux_x24_demux_io_out_1_bits_5; // @[Demux.scala 56:10]
  assign alu_io_input_bits_6 = accOutputDemux_x24_demux_io_out_1_bits_6; // @[Demux.scala 56:10]
  assign alu_io_input_bits_7 = accOutputDemux_x24_demux_io_out_1_bits_7; // @[Demux.scala 56:10]
  assign alu_io_input_bits_8 = accOutputDemux_x24_demux_io_out_1_bits_8; // @[Demux.scala 56:10]
  assign alu_io_input_bits_9 = accOutputDemux_x24_demux_io_out_1_bits_9; // @[Demux.scala 56:10]
  assign alu_io_input_bits_10 = accOutputDemux_x24_demux_io_out_1_bits_10; // @[Demux.scala 56:10]
  assign alu_io_input_bits_11 = accOutputDemux_x24_demux_io_out_1_bits_11; // @[Demux.scala 56:10]
  assign alu_io_input_bits_12 = accOutputDemux_x24_demux_io_out_1_bits_12; // @[Demux.scala 56:10]
  assign alu_io_input_bits_13 = accOutputDemux_x24_demux_io_out_1_bits_13; // @[Demux.scala 56:10]
  assign alu_io_input_bits_14 = accOutputDemux_x24_demux_io_out_1_bits_14; // @[Demux.scala 56:10]
  assign alu_io_input_bits_15 = accOutputDemux_x24_demux_io_out_1_bits_15; // @[Demux.scala 56:10]
  assign alu_io_input_bits_16 = accOutputDemux_x24_demux_io_out_1_bits_16; // @[Demux.scala 56:10]
  assign alu_io_input_bits_17 = accOutputDemux_x24_demux_io_out_1_bits_17; // @[Demux.scala 56:10]
  assign alu_io_input_bits_18 = accOutputDemux_x24_demux_io_out_1_bits_18; // @[Demux.scala 56:10]
  assign alu_io_input_bits_19 = accOutputDemux_x24_demux_io_out_1_bits_19; // @[Demux.scala 56:10]
  assign alu_io_input_bits_20 = accOutputDemux_x24_demux_io_out_1_bits_20; // @[Demux.scala 56:10]
  assign alu_io_input_bits_21 = accOutputDemux_x24_demux_io_out_1_bits_21; // @[Demux.scala 56:10]
  assign alu_io_input_bits_22 = accOutputDemux_x24_demux_io_out_1_bits_22; // @[Demux.scala 56:10]
  assign alu_io_input_bits_23 = accOutputDemux_x24_demux_io_out_1_bits_23; // @[Demux.scala 56:10]
  assign alu_io_input_bits_24 = accOutputDemux_x24_demux_io_out_1_bits_24; // @[Demux.scala 56:10]
  assign alu_io_input_bits_25 = accOutputDemux_x24_demux_io_out_1_bits_25; // @[Demux.scala 56:10]
  assign alu_io_input_bits_26 = accOutputDemux_x24_demux_io_out_1_bits_26; // @[Demux.scala 56:10]
  assign alu_io_input_bits_27 = accOutputDemux_x24_demux_io_out_1_bits_27; // @[Demux.scala 56:10]
  assign alu_io_input_bits_28 = accOutputDemux_x24_demux_io_out_1_bits_28; // @[Demux.scala 56:10]
  assign alu_io_input_bits_29 = accOutputDemux_x24_demux_io_out_1_bits_29; // @[Demux.scala 56:10]
  assign alu_io_input_bits_30 = accOutputDemux_x24_demux_io_out_1_bits_30; // @[Demux.scala 56:10]
  assign alu_io_input_bits_31 = accOutputDemux_x24_demux_io_out_1_bits_31; // @[Demux.scala 56:10]
  assign alu_io_output_ready = aluOutputDemux_x6_demux_io_in_ready; // @[Demux.scala 54:17]
  assign alu_io_instruction_valid = isNoOp ? 1'h0 : _GEN_169; // @[AccumulatorWithALUArray.scala 133:16 package.scala 405:15]
  assign alu_io_instruction_bits_op = isNoOp ? 4'h0 : _GEN_170; // @[AccumulatorWithALUArray.scala 133:16 package.scala 404:14]
  assign alu_io_instruction_bits_sourceLeft = isNoOp ? 1'h0 : _GEN_171; // @[AccumulatorWithALUArray.scala 133:16 package.scala 404:14]
  assign alu_io_instruction_bits_sourceRight = isNoOp ? 1'h0 : _GEN_172; // @[AccumulatorWithALUArray.scala 133:16 package.scala 404:14]
  assign alu_io_instruction_bits_dest = isNoOp ? 1'h0 : _GEN_173; // @[AccumulatorWithALUArray.scala 133:16 package.scala 404:14]
  assign aluOutputDemux_x6_demux_io_in_valid = alu_io_output_valid; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_0 = alu_io_output_bits_0; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_1 = alu_io_output_bits_1; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_2 = alu_io_output_bits_2; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_3 = alu_io_output_bits_3; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_4 = alu_io_output_bits_4; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_5 = alu_io_output_bits_5; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_6 = alu_io_output_bits_6; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_7 = alu_io_output_bits_7; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_8 = alu_io_output_bits_8; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_9 = alu_io_output_bits_9; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_10 = alu_io_output_bits_10; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_11 = alu_io_output_bits_11; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_12 = alu_io_output_bits_12; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_13 = alu_io_output_bits_13; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_14 = alu_io_output_bits_14; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_15 = alu_io_output_bits_15; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_16 = alu_io_output_bits_16; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_17 = alu_io_output_bits_17; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_18 = alu_io_output_bits_18; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_19 = alu_io_output_bits_19; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_20 = alu_io_output_bits_20; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_21 = alu_io_output_bits_21; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_22 = alu_io_output_bits_22; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_23 = alu_io_output_bits_23; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_24 = alu_io_output_bits_24; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_25 = alu_io_output_bits_25; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_26 = alu_io_output_bits_26; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_27 = alu_io_output_bits_27; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_28 = alu_io_output_bits_28; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_29 = alu_io_output_bits_29; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_30 = alu_io_output_bits_30; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_in_bits_31 = alu_io_output_bits_31; // @[Demux.scala 54:17]
  assign aluOutputDemux_x6_demux_io_sel_valid = aluOutputDemux_io_deq_valid; // @[Mem.scala 23:7]
  assign aluOutputDemux_x6_demux_io_sel_bits = aluOutputDemux_io_deq_bits; // @[Mem.scala 23:7]
  assign aluOutputDemux_x6_demux_io_out_0_ready = 1'h1; // @[Demux.scala 55:10]
  assign aluOutputDemux_x6_demux_io_out_1_ready = accInputMux_x15_mux_io_in_1_ready; // @[AccumulatorWithALUArray.scala 50:34 Mux.scala 80:18]
  assign aluOutputDemux_clock = clock;
  assign aluOutputDemux_reset = reset;
  assign aluOutputDemux_io_enq_valid = isNoOp ? 1'h0 : _GEN_156; // @[AccumulatorWithALUArray.scala 133:16 package.scala 405:15]
  assign aluOutputDemux_io_enq_bits = isNoOp ? 1'h0 : _GEN_48; // @[AccumulatorWithALUArray.scala 133:16 package.scala 404:14]
  assign aluOutputDemux_io_deq_ready = aluOutputDemux_x6_demux_io_sel_ready; // @[Mem.scala 23:7]
  assign accInputMux_x15_mux_io_in_0_valid = io_input_valid; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_0 = io_input_bits_0; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_1 = io_input_bits_1; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_2 = io_input_bits_2; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_3 = io_input_bits_3; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_4 = io_input_bits_4; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_5 = io_input_bits_5; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_6 = io_input_bits_6; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_7 = io_input_bits_7; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_8 = io_input_bits_8; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_9 = io_input_bits_9; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_10 = io_input_bits_10; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_11 = io_input_bits_11; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_12 = io_input_bits_12; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_13 = io_input_bits_13; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_14 = io_input_bits_14; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_15 = io_input_bits_15; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_16 = io_input_bits_16; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_17 = io_input_bits_17; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_18 = io_input_bits_18; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_19 = io_input_bits_19; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_20 = io_input_bits_20; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_21 = io_input_bits_21; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_22 = io_input_bits_22; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_23 = io_input_bits_23; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_24 = io_input_bits_24; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_25 = io_input_bits_25; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_26 = io_input_bits_26; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_27 = io_input_bits_27; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_28 = io_input_bits_28; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_29 = io_input_bits_29; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_30 = io_input_bits_30; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_0_bits_31 = io_input_bits_31; // @[Mux.scala 79:18]
  assign accInputMux_x15_mux_io_in_1_valid = aluOutputDemux_x6_demux_io_out_1_valid; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_0 = aluOutputDemux_x6_demux_io_out_1_bits_0; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_1 = aluOutputDemux_x6_demux_io_out_1_bits_1; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_2 = aluOutputDemux_x6_demux_io_out_1_bits_2; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_3 = aluOutputDemux_x6_demux_io_out_1_bits_3; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_4 = aluOutputDemux_x6_demux_io_out_1_bits_4; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_5 = aluOutputDemux_x6_demux_io_out_1_bits_5; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_6 = aluOutputDemux_x6_demux_io_out_1_bits_6; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_7 = aluOutputDemux_x6_demux_io_out_1_bits_7; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_8 = aluOutputDemux_x6_demux_io_out_1_bits_8; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_9 = aluOutputDemux_x6_demux_io_out_1_bits_9; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_10 = aluOutputDemux_x6_demux_io_out_1_bits_10; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_11 = aluOutputDemux_x6_demux_io_out_1_bits_11; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_12 = aluOutputDemux_x6_demux_io_out_1_bits_12; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_13 = aluOutputDemux_x6_demux_io_out_1_bits_13; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_14 = aluOutputDemux_x6_demux_io_out_1_bits_14; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_15 = aluOutputDemux_x6_demux_io_out_1_bits_15; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_16 = aluOutputDemux_x6_demux_io_out_1_bits_16; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_17 = aluOutputDemux_x6_demux_io_out_1_bits_17; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_18 = aluOutputDemux_x6_demux_io_out_1_bits_18; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_19 = aluOutputDemux_x6_demux_io_out_1_bits_19; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_20 = aluOutputDemux_x6_demux_io_out_1_bits_20; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_21 = aluOutputDemux_x6_demux_io_out_1_bits_21; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_22 = aluOutputDemux_x6_demux_io_out_1_bits_22; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_23 = aluOutputDemux_x6_demux_io_out_1_bits_23; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_24 = aluOutputDemux_x6_demux_io_out_1_bits_24; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_25 = aluOutputDemux_x6_demux_io_out_1_bits_25; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_26 = aluOutputDemux_x6_demux_io_out_1_bits_26; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_27 = aluOutputDemux_x6_demux_io_out_1_bits_27; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_28 = aluOutputDemux_x6_demux_io_out_1_bits_28; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_29 = aluOutputDemux_x6_demux_io_out_1_bits_29; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_30 = aluOutputDemux_x6_demux_io_out_1_bits_30; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_in_1_bits_31 = aluOutputDemux_x6_demux_io_out_1_bits_31; // @[AccumulatorWithALUArray.scala 50:34 Demux.scala 56:10]
  assign accInputMux_x15_mux_io_sel_valid = accInputMux_io_deq_valid; // @[Mem.scala 23:7]
  assign accInputMux_x15_mux_io_sel_bits = accInputMux_io_deq_bits; // @[Mem.scala 23:7]
  assign accInputMux_x15_mux_io_out_ready = acc_io_input_ready; // @[Mux.scala 81:9]
  assign accInputMux_clock = clock;
  assign accInputMux_reset = reset;
  assign accInputMux_io_enq_valid = isNoOp ? _GEN_50 : _GEN_159; // @[AccumulatorWithALUArray.scala 133:16]
  assign accInputMux_io_enq_bits = isNoOp ? 1'h0 : _GEN_48; // @[AccumulatorWithALUArray.scala 133:16]
  assign accInputMux_io_deq_ready = accInputMux_x15_mux_io_sel_ready; // @[Mem.scala 23:7]
  assign accOutputDemux_x24_demux_io_in_valid = acc_io_output_valid; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_0 = acc_io_output_bits_0; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_1 = acc_io_output_bits_1; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_2 = acc_io_output_bits_2; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_3 = acc_io_output_bits_3; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_4 = acc_io_output_bits_4; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_5 = acc_io_output_bits_5; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_6 = acc_io_output_bits_6; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_7 = acc_io_output_bits_7; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_8 = acc_io_output_bits_8; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_9 = acc_io_output_bits_9; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_10 = acc_io_output_bits_10; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_11 = acc_io_output_bits_11; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_12 = acc_io_output_bits_12; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_13 = acc_io_output_bits_13; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_14 = acc_io_output_bits_14; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_15 = acc_io_output_bits_15; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_16 = acc_io_output_bits_16; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_17 = acc_io_output_bits_17; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_18 = acc_io_output_bits_18; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_19 = acc_io_output_bits_19; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_20 = acc_io_output_bits_20; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_21 = acc_io_output_bits_21; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_22 = acc_io_output_bits_22; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_23 = acc_io_output_bits_23; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_24 = acc_io_output_bits_24; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_25 = acc_io_output_bits_25; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_26 = acc_io_output_bits_26; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_27 = acc_io_output_bits_27; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_28 = acc_io_output_bits_28; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_29 = acc_io_output_bits_29; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_30 = acc_io_output_bits_30; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_in_bits_31 = acc_io_output_bits_31; // @[Demux.scala 54:17]
  assign accOutputDemux_x24_demux_io_sel_valid = accOutputDemux_io_deq_valid; // @[Mem.scala 23:7]
  assign accOutputDemux_x24_demux_io_sel_bits = accOutputDemux_io_deq_bits; // @[Mem.scala 23:7]
  assign accOutputDemux_x24_demux_io_out_0_ready = io_output_ready; // @[Demux.scala 55:10]
  assign accOutputDemux_x24_demux_io_out_1_ready = alu_io_input_ready; // @[Demux.scala 56:10]
  assign accOutputDemux_clock = clock;
  assign accOutputDemux_reset = reset;
  assign accOutputDemux_io_enq_valid = isNoOp ? _GEN_57 : _GEN_166; // @[AccumulatorWithALUArray.scala 133:16]
  assign accOutputDemux_io_enq_bits = isNoOp ? 1'h0 : _GEN_167; // @[AccumulatorWithALUArray.scala 133:16]
  assign accOutputDemux_io_deq_ready = accOutputDemux_x24_demux_io_sel_ready; // @[Mem.scala 23:7]
  assign accWriteEnqueuer_clock = clock;
  assign accWriteEnqueuer_reset = reset;
  assign accWriteEnqueuer_io_in_valid = isNoOp & _GEN_43; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 40:17]
  assign accWriteEnqueuer_io_out_0_ready = isNoOp & _GEN_44; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign accWriteEnqueuer_io_out_1_ready = isNoOp & _GEN_49; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign accReadEnqueuer_clock = clock;
  assign accReadEnqueuer_reset = reset;
  assign accReadEnqueuer_io_in_valid = isNoOp & _GEN_54; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 40:17]
  assign accReadEnqueuer_io_out_0_ready = isNoOp & _GEN_55; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign accReadEnqueuer_io_out_1_ready = isNoOp & _GEN_56; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdRWWriteEnqueuer_clock = clock;
  assign simdRWWriteEnqueuer_reset = reset;
  assign simdRWWriteEnqueuer_io_in_valid = isNoOp ? 1'h0 : _GEN_149; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 40:17]
  assign simdRWWriteEnqueuer_io_out_0_ready = isNoOp ? 1'h0 : _GEN_150; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdRWWriteEnqueuer_io_out_1_ready = isNoOp ? 1'h0 : _GEN_155; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdRWWriteEnqueuer_io_out_2_ready = isNoOp ? 1'h0 : _GEN_158; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdRWReadEnqueuer_clock = clock;
  assign simdRWReadEnqueuer_reset = reset;
  assign simdRWReadEnqueuer_io_in_valid = isNoOp ? 1'h0 : _GEN_163; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 40:17]
  assign simdRWReadEnqueuer_io_out_0_ready = isNoOp ? 1'h0 : _GEN_164; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdRWReadEnqueuer_io_out_1_ready = isNoOp ? 1'h0 : _GEN_165; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdRWReadEnqueuer_io_out_2_ready = isNoOp ? 1'h0 : _GEN_168; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdWriteEnqueuer_clock = clock;
  assign simdWriteEnqueuer_reset = reset;
  assign simdWriteEnqueuer_io_in_valid = isNoOp ? 1'h0 : _GEN_179; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 40:17]
  assign simdWriteEnqueuer_io_out_0_ready = isNoOp ? 1'h0 : _GEN_180; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdWriteEnqueuer_io_out_1_ready = isNoOp ? 1'h0 : _GEN_181; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdWriteEnqueuer_io_out_2_ready = isNoOp ? 1'h0 : _GEN_182; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdWriteEnqueuer_io_out_3_ready = isNoOp ? 1'h0 : _GEN_183; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdReadEnqueuer_clock = clock;
  assign simdReadEnqueuer_reset = reset;
  assign simdReadEnqueuer_io_in_valid = isNoOp ? 1'h0 : _GEN_174; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 40:17]
  assign simdReadEnqueuer_io_out_0_ready = isNoOp ? 1'h0 : _GEN_175; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdReadEnqueuer_io_out_1_ready = isNoOp ? 1'h0 : _GEN_176; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdReadEnqueuer_io_out_2_ready = isNoOp ? 1'h0 : _GEN_177; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdReadEnqueuer_io_out_3_ready = isNoOp ? 1'h0 : _GEN_178; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdEnqueuer_clock = clock;
  assign simdEnqueuer_reset = reset;
  assign simdEnqueuer_io_in_valid = isNoOp ? 1'h0 : _GEN_184; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 40:17]
  assign simdEnqueuer_io_out_0_ready = isNoOp ? 1'h0 : _GEN_185; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  assign simdEnqueuer_io_out_1_ready = isNoOp ? 1'h0 : _GEN_186; // @[AccumulatorWithALUArray.scala 133:16 MultiEnqueue.scala 42:18]
  always @(posedge clock) begin
    if (reset) begin // @[AccumulatorWithALUArray.scala 110:29]
      readEnqueued <= 1'h0; // @[AccumulatorWithALUArray.scala 110:29]
    end else if (isNoOp) begin // @[AccumulatorWithALUArray.scala 133:16]
      readEnqueued <= _GEN_53;
    end else begin
      readEnqueued <= _GEN_162;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  readEnqueued = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InnerDualPortMem_1(
  input         clock,
  input         reset,
  input  [13:0] io_portA_address,
  input         io_portA_read_enable,
  output [15:0] io_portA_read_data_0,
  output [15:0] io_portA_read_data_1,
  output [15:0] io_portA_read_data_2,
  output [15:0] io_portA_read_data_3,
  output [15:0] io_portA_read_data_4,
  output [15:0] io_portA_read_data_5,
  output [15:0] io_portA_read_data_6,
  output [15:0] io_portA_read_data_7,
  output [15:0] io_portA_read_data_8,
  output [15:0] io_portA_read_data_9,
  output [15:0] io_portA_read_data_10,
  output [15:0] io_portA_read_data_11,
  output [15:0] io_portA_read_data_12,
  output [15:0] io_portA_read_data_13,
  output [15:0] io_portA_read_data_14,
  output [15:0] io_portA_read_data_15,
  output [15:0] io_portA_read_data_16,
  output [15:0] io_portA_read_data_17,
  output [15:0] io_portA_read_data_18,
  output [15:0] io_portA_read_data_19,
  output [15:0] io_portA_read_data_20,
  output [15:0] io_portA_read_data_21,
  output [15:0] io_portA_read_data_22,
  output [15:0] io_portA_read_data_23,
  output [15:0] io_portA_read_data_24,
  output [15:0] io_portA_read_data_25,
  output [15:0] io_portA_read_data_26,
  output [15:0] io_portA_read_data_27,
  output [15:0] io_portA_read_data_28,
  output [15:0] io_portA_read_data_29,
  output [15:0] io_portA_read_data_30,
  output [15:0] io_portA_read_data_31,
  input         io_portA_write_enable,
  input  [15:0] io_portA_write_data_0,
  input  [15:0] io_portA_write_data_1,
  input  [15:0] io_portA_write_data_2,
  input  [15:0] io_portA_write_data_3,
  input  [15:0] io_portA_write_data_4,
  input  [15:0] io_portA_write_data_5,
  input  [15:0] io_portA_write_data_6,
  input  [15:0] io_portA_write_data_7,
  input  [15:0] io_portA_write_data_8,
  input  [15:0] io_portA_write_data_9,
  input  [15:0] io_portA_write_data_10,
  input  [15:0] io_portA_write_data_11,
  input  [15:0] io_portA_write_data_12,
  input  [15:0] io_portA_write_data_13,
  input  [15:0] io_portA_write_data_14,
  input  [15:0] io_portA_write_data_15,
  input  [15:0] io_portA_write_data_16,
  input  [15:0] io_portA_write_data_17,
  input  [15:0] io_portA_write_data_18,
  input  [15:0] io_portA_write_data_19,
  input  [15:0] io_portA_write_data_20,
  input  [15:0] io_portA_write_data_21,
  input  [15:0] io_portA_write_data_22,
  input  [15:0] io_portA_write_data_23,
  input  [15:0] io_portA_write_data_24,
  input  [15:0] io_portA_write_data_25,
  input  [15:0] io_portA_write_data_26,
  input  [15:0] io_portA_write_data_27,
  input  [15:0] io_portA_write_data_28,
  input  [15:0] io_portA_write_data_29,
  input  [15:0] io_portA_write_data_30,
  input  [15:0] io_portA_write_data_31,
  input  [13:0] io_portB_address,
  input         io_portB_read_enable,
  output [15:0] io_portB_read_data_0,
  output [15:0] io_portB_read_data_1,
  output [15:0] io_portB_read_data_2,
  output [15:0] io_portB_read_data_3,
  output [15:0] io_portB_read_data_4,
  output [15:0] io_portB_read_data_5,
  output [15:0] io_portB_read_data_6,
  output [15:0] io_portB_read_data_7,
  output [15:0] io_portB_read_data_8,
  output [15:0] io_portB_read_data_9,
  output [15:0] io_portB_read_data_10,
  output [15:0] io_portB_read_data_11,
  output [15:0] io_portB_read_data_12,
  output [15:0] io_portB_read_data_13,
  output [15:0] io_portB_read_data_14,
  output [15:0] io_portB_read_data_15,
  output [15:0] io_portB_read_data_16,
  output [15:0] io_portB_read_data_17,
  output [15:0] io_portB_read_data_18,
  output [15:0] io_portB_read_data_19,
  output [15:0] io_portB_read_data_20,
  output [15:0] io_portB_read_data_21,
  output [15:0] io_portB_read_data_22,
  output [15:0] io_portB_read_data_23,
  output [15:0] io_portB_read_data_24,
  output [15:0] io_portB_read_data_25,
  output [15:0] io_portB_read_data_26,
  output [15:0] io_portB_read_data_27,
  output [15:0] io_portB_read_data_28,
  output [15:0] io_portB_read_data_29,
  output [15:0] io_portB_read_data_30,
  output [15:0] io_portB_read_data_31,
  input         io_portB_write_enable,
  input  [15:0] io_portB_write_data_0,
  input  [15:0] io_portB_write_data_1,
  input  [15:0] io_portB_write_data_2,
  input  [15:0] io_portB_write_data_3,
  input  [15:0] io_portB_write_data_4,
  input  [15:0] io_portB_write_data_5,
  input  [15:0] io_portB_write_data_6,
  input  [15:0] io_portB_write_data_7,
  input  [15:0] io_portB_write_data_8,
  input  [15:0] io_portB_write_data_9,
  input  [15:0] io_portB_write_data_10,
  input  [15:0] io_portB_write_data_11,
  input  [15:0] io_portB_write_data_12,
  input  [15:0] io_portB_write_data_13,
  input  [15:0] io_portB_write_data_14,
  input  [15:0] io_portB_write_data_15,
  input  [15:0] io_portB_write_data_16,
  input  [15:0] io_portB_write_data_17,
  input  [15:0] io_portB_write_data_18,
  input  [15:0] io_portB_write_data_19,
  input  [15:0] io_portB_write_data_20,
  input  [15:0] io_portB_write_data_21,
  input  [15:0] io_portB_write_data_22,
  input  [15:0] io_portB_write_data_23,
  input  [15:0] io_portB_write_data_24,
  input  [15:0] io_portB_write_data_25,
  input  [15:0] io_portB_write_data_26,
  input  [15:0] io_portB_write_data_27,
  input  [15:0] io_portB_write_data_28,
  input  [15:0] io_portB_write_data_29,
  input  [15:0] io_portB_write_data_30,
  input  [15:0] io_portB_write_data_31
);
  wire  mem_clka; // @[DualPortMem.scala 173:25]
  wire  mem_wea; // @[DualPortMem.scala 173:25]
  wire  mem_ena; // @[DualPortMem.scala 173:25]
  wire [13:0] mem_addra; // @[DualPortMem.scala 173:25]
  wire [511:0] mem_dia; // @[DualPortMem.scala 173:25]
  wire [511:0] mem_doa; // @[DualPortMem.scala 173:25]
  wire  mem_clkb; // @[DualPortMem.scala 173:25]
  wire  mem_web; // @[DualPortMem.scala 173:25]
  wire  mem_enb; // @[DualPortMem.scala 173:25]
  wire [13:0] mem_addrb; // @[DualPortMem.scala 173:25]
  wire [511:0] mem_dib; // @[DualPortMem.scala 173:25]
  wire [511:0] mem_dob; // @[DualPortMem.scala 173:25]
  wire [511:0] _io_portA_read_data_WIRE_1 = mem_doa;
  wire [127:0] mem_io_dia_lo_lo = {io_portA_write_data_7,io_portA_write_data_6,io_portA_write_data_5,
    io_portA_write_data_4,io_portA_write_data_3,io_portA_write_data_2,io_portA_write_data_1,io_portA_write_data_0}; // @[DualPortMem.scala 180:51]
  wire [255:0] mem_io_dia_lo = {io_portA_write_data_15,io_portA_write_data_14,io_portA_write_data_13,
    io_portA_write_data_12,io_portA_write_data_11,io_portA_write_data_10,io_portA_write_data_9,io_portA_write_data_8,
    mem_io_dia_lo_lo}; // @[DualPortMem.scala 180:51]
  wire [127:0] mem_io_dia_hi_lo = {io_portA_write_data_23,io_portA_write_data_22,io_portA_write_data_21,
    io_portA_write_data_20,io_portA_write_data_19,io_portA_write_data_18,io_portA_write_data_17,io_portA_write_data_16}; // @[DualPortMem.scala 180:51]
  wire [255:0] mem_io_dia_hi = {io_portA_write_data_31,io_portA_write_data_30,io_portA_write_data_29,
    io_portA_write_data_28,io_portA_write_data_27,io_portA_write_data_26,io_portA_write_data_25,io_portA_write_data_24,
    mem_io_dia_hi_lo}; // @[DualPortMem.scala 180:51]
  wire [511:0] _io_portB_read_data_WIRE_1 = mem_dob;
  wire [127:0] mem_io_dib_lo_lo = {io_portB_write_data_7,io_portB_write_data_6,io_portB_write_data_5,
    io_portB_write_data_4,io_portB_write_data_3,io_portB_write_data_2,io_portB_write_data_1,io_portB_write_data_0}; // @[DualPortMem.scala 187:51]
  wire [255:0] mem_io_dib_lo = {io_portB_write_data_15,io_portB_write_data_14,io_portB_write_data_13,
    io_portB_write_data_12,io_portB_write_data_11,io_portB_write_data_10,io_portB_write_data_9,io_portB_write_data_8,
    mem_io_dib_lo_lo}; // @[DualPortMem.scala 187:51]
  wire [127:0] mem_io_dib_hi_lo = {io_portB_write_data_23,io_portB_write_data_22,io_portB_write_data_21,
    io_portB_write_data_20,io_portB_write_data_19,io_portB_write_data_18,io_portB_write_data_17,io_portB_write_data_16}; // @[DualPortMem.scala 187:51]
  wire [255:0] mem_io_dib_hi = {io_portB_write_data_31,io_portB_write_data_30,io_portB_write_data_29,
    io_portB_write_data_28,io_portB_write_data_27,io_portB_write_data_26,io_portB_write_data_25,io_portB_write_data_24,
    mem_io_dib_hi_lo}; // @[DualPortMem.scala 187:51]
  bram_dp_512x16384 mem ( // @[DualPortMem.scala 173:25]
    .clka(mem_clka),
    .wea(mem_wea),
    .ena(mem_ena),
    .addra(mem_addra),
    .dia(mem_dia),
    .doa(mem_doa),
    .clkb(mem_clkb),
    .web(mem_web),
    .enb(mem_enb),
    .addrb(mem_addrb),
    .dib(mem_dib),
    .dob(mem_dob)
  );
  assign io_portA_read_data_0 = _io_portA_read_data_WIRE_1[15:0]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_1 = _io_portA_read_data_WIRE_1[31:16]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_2 = _io_portA_read_data_WIRE_1[47:32]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_3 = _io_portA_read_data_WIRE_1[63:48]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_4 = _io_portA_read_data_WIRE_1[79:64]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_5 = _io_portA_read_data_WIRE_1[95:80]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_6 = _io_portA_read_data_WIRE_1[111:96]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_7 = _io_portA_read_data_WIRE_1[127:112]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_8 = _io_portA_read_data_WIRE_1[143:128]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_9 = _io_portA_read_data_WIRE_1[159:144]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_10 = _io_portA_read_data_WIRE_1[175:160]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_11 = _io_portA_read_data_WIRE_1[191:176]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_12 = _io_portA_read_data_WIRE_1[207:192]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_13 = _io_portA_read_data_WIRE_1[223:208]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_14 = _io_portA_read_data_WIRE_1[239:224]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_15 = _io_portA_read_data_WIRE_1[255:240]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_16 = _io_portA_read_data_WIRE_1[271:256]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_17 = _io_portA_read_data_WIRE_1[287:272]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_18 = _io_portA_read_data_WIRE_1[303:288]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_19 = _io_portA_read_data_WIRE_1[319:304]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_20 = _io_portA_read_data_WIRE_1[335:320]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_21 = _io_portA_read_data_WIRE_1[351:336]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_22 = _io_portA_read_data_WIRE_1[367:352]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_23 = _io_portA_read_data_WIRE_1[383:368]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_24 = _io_portA_read_data_WIRE_1[399:384]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_25 = _io_portA_read_data_WIRE_1[415:400]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_26 = _io_portA_read_data_WIRE_1[431:416]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_27 = _io_portA_read_data_WIRE_1[447:432]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_28 = _io_portA_read_data_WIRE_1[463:448]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_29 = _io_portA_read_data_WIRE_1[479:464]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_30 = _io_portA_read_data_WIRE_1[495:480]; // @[DualPortMem.scala 178:50]
  assign io_portA_read_data_31 = _io_portA_read_data_WIRE_1[511:496]; // @[DualPortMem.scala 178:50]
  assign io_portB_read_data_0 = _io_portB_read_data_WIRE_1[15:0]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_1 = _io_portB_read_data_WIRE_1[31:16]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_2 = _io_portB_read_data_WIRE_1[47:32]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_3 = _io_portB_read_data_WIRE_1[63:48]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_4 = _io_portB_read_data_WIRE_1[79:64]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_5 = _io_portB_read_data_WIRE_1[95:80]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_6 = _io_portB_read_data_WIRE_1[111:96]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_7 = _io_portB_read_data_WIRE_1[127:112]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_8 = _io_portB_read_data_WIRE_1[143:128]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_9 = _io_portB_read_data_WIRE_1[159:144]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_10 = _io_portB_read_data_WIRE_1[175:160]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_11 = _io_portB_read_data_WIRE_1[191:176]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_12 = _io_portB_read_data_WIRE_1[207:192]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_13 = _io_portB_read_data_WIRE_1[223:208]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_14 = _io_portB_read_data_WIRE_1[239:224]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_15 = _io_portB_read_data_WIRE_1[255:240]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_16 = _io_portB_read_data_WIRE_1[271:256]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_17 = _io_portB_read_data_WIRE_1[287:272]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_18 = _io_portB_read_data_WIRE_1[303:288]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_19 = _io_portB_read_data_WIRE_1[319:304]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_20 = _io_portB_read_data_WIRE_1[335:320]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_21 = _io_portB_read_data_WIRE_1[351:336]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_22 = _io_portB_read_data_WIRE_1[367:352]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_23 = _io_portB_read_data_WIRE_1[383:368]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_24 = _io_portB_read_data_WIRE_1[399:384]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_25 = _io_portB_read_data_WIRE_1[415:400]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_26 = _io_portB_read_data_WIRE_1[431:416]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_27 = _io_portB_read_data_WIRE_1[447:432]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_28 = _io_portB_read_data_WIRE_1[463:448]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_29 = _io_portB_read_data_WIRE_1[479:464]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_30 = _io_portB_read_data_WIRE_1[495:480]; // @[DualPortMem.scala 185:50]
  assign io_portB_read_data_31 = _io_portB_read_data_WIRE_1[511:496]; // @[DualPortMem.scala 185:50]
  assign mem_clka = clock; // @[DualPortMem.scala 175:30]
  assign mem_wea = io_portA_write_enable; // @[DualPortMem.scala 179:20]
  assign mem_ena = ~reset; // @[DualPortMem.scala 176:23]
  assign mem_addra = io_portA_address; // @[DualPortMem.scala 177:22]
  assign mem_dia = {mem_io_dia_hi,mem_io_dia_lo}; // @[DualPortMem.scala 180:51]
  assign mem_clkb = clock; // @[DualPortMem.scala 182:30]
  assign mem_web = io_portB_write_enable; // @[DualPortMem.scala 186:20]
  assign mem_enb = ~reset; // @[DualPortMem.scala 183:23]
  assign mem_addrb = io_portB_address; // @[DualPortMem.scala 184:22]
  assign mem_dib = {mem_io_dib_hi,mem_io_dib_lo}; // @[DualPortMem.scala 187:51]
endmodule
module DualPortMem_1(
  input         clock,
  input         reset,
  output        io_portA_control_ready,
  input         io_portA_control_valid,
  input         io_portA_control_bits_write,
  input  [13:0] io_portA_control_bits_address,
  output        io_portA_input_ready,
  input         io_portA_input_valid,
  input  [15:0] io_portA_input_bits_0,
  input  [15:0] io_portA_input_bits_1,
  input  [15:0] io_portA_input_bits_2,
  input  [15:0] io_portA_input_bits_3,
  input  [15:0] io_portA_input_bits_4,
  input  [15:0] io_portA_input_bits_5,
  input  [15:0] io_portA_input_bits_6,
  input  [15:0] io_portA_input_bits_7,
  input  [15:0] io_portA_input_bits_8,
  input  [15:0] io_portA_input_bits_9,
  input  [15:0] io_portA_input_bits_10,
  input  [15:0] io_portA_input_bits_11,
  input  [15:0] io_portA_input_bits_12,
  input  [15:0] io_portA_input_bits_13,
  input  [15:0] io_portA_input_bits_14,
  input  [15:0] io_portA_input_bits_15,
  input  [15:0] io_portA_input_bits_16,
  input  [15:0] io_portA_input_bits_17,
  input  [15:0] io_portA_input_bits_18,
  input  [15:0] io_portA_input_bits_19,
  input  [15:0] io_portA_input_bits_20,
  input  [15:0] io_portA_input_bits_21,
  input  [15:0] io_portA_input_bits_22,
  input  [15:0] io_portA_input_bits_23,
  input  [15:0] io_portA_input_bits_24,
  input  [15:0] io_portA_input_bits_25,
  input  [15:0] io_portA_input_bits_26,
  input  [15:0] io_portA_input_bits_27,
  input  [15:0] io_portA_input_bits_28,
  input  [15:0] io_portA_input_bits_29,
  input  [15:0] io_portA_input_bits_30,
  input  [15:0] io_portA_input_bits_31,
  input         io_portA_output_ready,
  output        io_portA_output_valid,
  output [15:0] io_portA_output_bits_0,
  output [15:0] io_portA_output_bits_1,
  output [15:0] io_portA_output_bits_2,
  output [15:0] io_portA_output_bits_3,
  output [15:0] io_portA_output_bits_4,
  output [15:0] io_portA_output_bits_5,
  output [15:0] io_portA_output_bits_6,
  output [15:0] io_portA_output_bits_7,
  output [15:0] io_portA_output_bits_8,
  output [15:0] io_portA_output_bits_9,
  output [15:0] io_portA_output_bits_10,
  output [15:0] io_portA_output_bits_11,
  output [15:0] io_portA_output_bits_12,
  output [15:0] io_portA_output_bits_13,
  output [15:0] io_portA_output_bits_14,
  output [15:0] io_portA_output_bits_15,
  output [15:0] io_portA_output_bits_16,
  output [15:0] io_portA_output_bits_17,
  output [15:0] io_portA_output_bits_18,
  output [15:0] io_portA_output_bits_19,
  output [15:0] io_portA_output_bits_20,
  output [15:0] io_portA_output_bits_21,
  output [15:0] io_portA_output_bits_22,
  output [15:0] io_portA_output_bits_23,
  output [15:0] io_portA_output_bits_24,
  output [15:0] io_portA_output_bits_25,
  output [15:0] io_portA_output_bits_26,
  output [15:0] io_portA_output_bits_27,
  output [15:0] io_portA_output_bits_28,
  output [15:0] io_portA_output_bits_29,
  output [15:0] io_portA_output_bits_30,
  output [15:0] io_portA_output_bits_31,
  output        io_portB_control_ready,
  input         io_portB_control_valid,
  input         io_portB_control_bits_write,
  input  [13:0] io_portB_control_bits_address,
  output        io_portB_input_ready,
  input         io_portB_input_valid,
  input  [15:0] io_portB_input_bits_0,
  input  [15:0] io_portB_input_bits_1,
  input  [15:0] io_portB_input_bits_2,
  input  [15:0] io_portB_input_bits_3,
  input  [15:0] io_portB_input_bits_4,
  input  [15:0] io_portB_input_bits_5,
  input  [15:0] io_portB_input_bits_6,
  input  [15:0] io_portB_input_bits_7,
  input  [15:0] io_portB_input_bits_8,
  input  [15:0] io_portB_input_bits_9,
  input  [15:0] io_portB_input_bits_10,
  input  [15:0] io_portB_input_bits_11,
  input  [15:0] io_portB_input_bits_12,
  input  [15:0] io_portB_input_bits_13,
  input  [15:0] io_portB_input_bits_14,
  input  [15:0] io_portB_input_bits_15,
  input  [15:0] io_portB_input_bits_16,
  input  [15:0] io_portB_input_bits_17,
  input  [15:0] io_portB_input_bits_18,
  input  [15:0] io_portB_input_bits_19,
  input  [15:0] io_portB_input_bits_20,
  input  [15:0] io_portB_input_bits_21,
  input  [15:0] io_portB_input_bits_22,
  input  [15:0] io_portB_input_bits_23,
  input  [15:0] io_portB_input_bits_24,
  input  [15:0] io_portB_input_bits_25,
  input  [15:0] io_portB_input_bits_26,
  input  [15:0] io_portB_input_bits_27,
  input  [15:0] io_portB_input_bits_28,
  input  [15:0] io_portB_input_bits_29,
  input  [15:0] io_portB_input_bits_30,
  input  [15:0] io_portB_input_bits_31,
  input         io_portB_output_ready,
  output        io_portB_output_valid,
  output [15:0] io_portB_output_bits_0,
  output [15:0] io_portB_output_bits_1,
  output [15:0] io_portB_output_bits_2,
  output [15:0] io_portB_output_bits_3,
  output [15:0] io_portB_output_bits_4,
  output [15:0] io_portB_output_bits_5,
  output [15:0] io_portB_output_bits_6,
  output [15:0] io_portB_output_bits_7,
  output [15:0] io_portB_output_bits_8,
  output [15:0] io_portB_output_bits_9,
  output [15:0] io_portB_output_bits_10,
  output [15:0] io_portB_output_bits_11,
  output [15:0] io_portB_output_bits_12,
  output [15:0] io_portB_output_bits_13,
  output [15:0] io_portB_output_bits_14,
  output [15:0] io_portB_output_bits_15,
  output [15:0] io_portB_output_bits_16,
  output [15:0] io_portB_output_bits_17,
  output [15:0] io_portB_output_bits_18,
  output [15:0] io_portB_output_bits_19,
  output [15:0] io_portB_output_bits_20,
  output [15:0] io_portB_output_bits_21,
  output [15:0] io_portB_output_bits_22,
  output [15:0] io_portB_output_bits_23,
  output [15:0] io_portB_output_bits_24,
  output [15:0] io_portB_output_bits_25,
  output [15:0] io_portB_output_bits_26,
  output [15:0] io_portB_output_bits_27,
  output [15:0] io_portB_output_bits_28,
  output [15:0] io_portB_output_bits_29,
  output [15:0] io_portB_output_bits_30,
  output [15:0] io_portB_output_bits_31,
  input         io_tracepoint,
  input  [31:0] io_programCounter
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  mem_clock; // @[DualPortMem.scala 33:19]
  wire  mem_reset; // @[DualPortMem.scala 33:19]
  wire [13:0] mem_io_portA_address; // @[DualPortMem.scala 33:19]
  wire  mem_io_portA_read_enable; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_0; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_1; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_2; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_3; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_4; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_5; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_6; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_7; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_8; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_9; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_10; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_11; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_12; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_13; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_14; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_15; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_16; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_17; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_18; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_19; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_20; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_21; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_22; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_23; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_24; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_25; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_26; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_27; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_28; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_29; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_30; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_read_data_31; // @[DualPortMem.scala 33:19]
  wire  mem_io_portA_write_enable; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_0; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_1; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_2; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_3; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_4; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_5; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_6; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_7; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_8; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_9; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_10; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_11; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_12; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_13; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_14; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_15; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_16; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_17; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_18; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_19; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_20; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_21; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_22; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_23; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_24; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_25; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_26; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_27; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_28; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_29; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_30; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portA_write_data_31; // @[DualPortMem.scala 33:19]
  wire [13:0] mem_io_portB_address; // @[DualPortMem.scala 33:19]
  wire  mem_io_portB_read_enable; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_0; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_1; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_2; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_3; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_4; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_5; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_6; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_7; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_8; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_9; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_10; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_11; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_12; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_13; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_14; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_15; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_16; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_17; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_18; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_19; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_20; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_21; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_22; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_23; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_24; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_25; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_26; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_27; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_28; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_29; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_30; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_read_data_31; // @[DualPortMem.scala 33:19]
  wire  mem_io_portB_write_enable; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_0; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_1; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_2; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_3; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_4; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_5; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_6; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_7; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_8; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_9; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_10; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_11; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_12; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_13; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_14; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_15; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_16; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_17; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_18; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_19; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_20; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_21; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_22; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_23; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_24; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_25; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_26; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_27; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_28; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_29; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_30; // @[DualPortMem.scala 33:19]
  wire [15:0] mem_io_portB_write_data_31; // @[DualPortMem.scala 33:19]
  wire  output__clock; // @[DualPortMem.scala 48:24]
  wire  output__reset; // @[DualPortMem.scala 48:24]
  wire  output__io_enq_ready; // @[DualPortMem.scala 48:24]
  wire  output__io_enq_valid; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_0; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_1; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_2; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_3; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_4; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_5; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_6; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_7; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_8; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_9; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_10; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_11; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_12; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_13; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_14; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_15; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_16; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_17; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_18; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_19; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_20; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_21; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_22; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_23; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_24; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_25; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_26; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_27; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_28; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_29; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_30; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_enq_bits_31; // @[DualPortMem.scala 48:24]
  wire  output__io_deq_ready; // @[DualPortMem.scala 48:24]
  wire  output__io_deq_valid; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_0; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_1; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_2; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_3; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_4; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_5; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_6; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_7; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_8; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_9; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_10; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_11; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_12; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_13; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_14; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_15; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_16; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_17; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_18; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_19; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_20; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_21; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_22; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_23; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_24; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_25; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_26; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_27; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_28; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_29; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_30; // @[DualPortMem.scala 48:24]
  wire [15:0] output__io_deq_bits_31; // @[DualPortMem.scala 48:24]
  wire [1:0] output__io_count; // @[DualPortMem.scala 48:24]
  wire  output_1_clock; // @[DualPortMem.scala 48:24]
  wire  output_1_reset; // @[DualPortMem.scala 48:24]
  wire  output_1_io_enq_ready; // @[DualPortMem.scala 48:24]
  wire  output_1_io_enq_valid; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_0; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_1; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_2; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_3; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_4; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_5; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_6; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_7; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_8; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_9; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_10; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_11; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_12; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_13; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_14; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_15; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_16; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_17; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_18; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_19; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_20; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_21; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_22; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_23; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_24; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_25; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_26; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_27; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_28; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_29; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_30; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_enq_bits_31; // @[DualPortMem.scala 48:24]
  wire  output_1_io_deq_ready; // @[DualPortMem.scala 48:24]
  wire  output_1_io_deq_valid; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_0; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_1; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_2; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_3; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_4; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_5; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_6; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_7; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_8; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_9; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_10; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_11; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_12; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_13; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_14; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_15; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_16; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_17; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_18; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_19; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_20; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_21; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_22; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_23; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_24; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_25; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_26; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_27; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_28; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_29; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_30; // @[DualPortMem.scala 48:24]
  wire [15:0] output_1_io_deq_bits_31; // @[DualPortMem.scala 48:24]
  wire [1:0] output_1_io_count; // @[DualPortMem.scala 48:24]
  wire  outputReady = output__io_count < 2'h2; // @[DualPortMem.scala 55:39]
  reg  output_io_enq_valid_sr_0; // @[ShiftRegister.scala 10:22]
  wire  outputReady_1 = output_1_io_count < 2'h2; // @[DualPortMem.scala 55:39]
  reg  output_io_enq_valid_sr_1_0; // @[ShiftRegister.scala 10:22]
  InnerDualPortMem_1 mem ( // @[DualPortMem.scala 33:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_portA_address(mem_io_portA_address),
    .io_portA_read_enable(mem_io_portA_read_enable),
    .io_portA_read_data_0(mem_io_portA_read_data_0),
    .io_portA_read_data_1(mem_io_portA_read_data_1),
    .io_portA_read_data_2(mem_io_portA_read_data_2),
    .io_portA_read_data_3(mem_io_portA_read_data_3),
    .io_portA_read_data_4(mem_io_portA_read_data_4),
    .io_portA_read_data_5(mem_io_portA_read_data_5),
    .io_portA_read_data_6(mem_io_portA_read_data_6),
    .io_portA_read_data_7(mem_io_portA_read_data_7),
    .io_portA_read_data_8(mem_io_portA_read_data_8),
    .io_portA_read_data_9(mem_io_portA_read_data_9),
    .io_portA_read_data_10(mem_io_portA_read_data_10),
    .io_portA_read_data_11(mem_io_portA_read_data_11),
    .io_portA_read_data_12(mem_io_portA_read_data_12),
    .io_portA_read_data_13(mem_io_portA_read_data_13),
    .io_portA_read_data_14(mem_io_portA_read_data_14),
    .io_portA_read_data_15(mem_io_portA_read_data_15),
    .io_portA_read_data_16(mem_io_portA_read_data_16),
    .io_portA_read_data_17(mem_io_portA_read_data_17),
    .io_portA_read_data_18(mem_io_portA_read_data_18),
    .io_portA_read_data_19(mem_io_portA_read_data_19),
    .io_portA_read_data_20(mem_io_portA_read_data_20),
    .io_portA_read_data_21(mem_io_portA_read_data_21),
    .io_portA_read_data_22(mem_io_portA_read_data_22),
    .io_portA_read_data_23(mem_io_portA_read_data_23),
    .io_portA_read_data_24(mem_io_portA_read_data_24),
    .io_portA_read_data_25(mem_io_portA_read_data_25),
    .io_portA_read_data_26(mem_io_portA_read_data_26),
    .io_portA_read_data_27(mem_io_portA_read_data_27),
    .io_portA_read_data_28(mem_io_portA_read_data_28),
    .io_portA_read_data_29(mem_io_portA_read_data_29),
    .io_portA_read_data_30(mem_io_portA_read_data_30),
    .io_portA_read_data_31(mem_io_portA_read_data_31),
    .io_portA_write_enable(mem_io_portA_write_enable),
    .io_portA_write_data_0(mem_io_portA_write_data_0),
    .io_portA_write_data_1(mem_io_portA_write_data_1),
    .io_portA_write_data_2(mem_io_portA_write_data_2),
    .io_portA_write_data_3(mem_io_portA_write_data_3),
    .io_portA_write_data_4(mem_io_portA_write_data_4),
    .io_portA_write_data_5(mem_io_portA_write_data_5),
    .io_portA_write_data_6(mem_io_portA_write_data_6),
    .io_portA_write_data_7(mem_io_portA_write_data_7),
    .io_portA_write_data_8(mem_io_portA_write_data_8),
    .io_portA_write_data_9(mem_io_portA_write_data_9),
    .io_portA_write_data_10(mem_io_portA_write_data_10),
    .io_portA_write_data_11(mem_io_portA_write_data_11),
    .io_portA_write_data_12(mem_io_portA_write_data_12),
    .io_portA_write_data_13(mem_io_portA_write_data_13),
    .io_portA_write_data_14(mem_io_portA_write_data_14),
    .io_portA_write_data_15(mem_io_portA_write_data_15),
    .io_portA_write_data_16(mem_io_portA_write_data_16),
    .io_portA_write_data_17(mem_io_portA_write_data_17),
    .io_portA_write_data_18(mem_io_portA_write_data_18),
    .io_portA_write_data_19(mem_io_portA_write_data_19),
    .io_portA_write_data_20(mem_io_portA_write_data_20),
    .io_portA_write_data_21(mem_io_portA_write_data_21),
    .io_portA_write_data_22(mem_io_portA_write_data_22),
    .io_portA_write_data_23(mem_io_portA_write_data_23),
    .io_portA_write_data_24(mem_io_portA_write_data_24),
    .io_portA_write_data_25(mem_io_portA_write_data_25),
    .io_portA_write_data_26(mem_io_portA_write_data_26),
    .io_portA_write_data_27(mem_io_portA_write_data_27),
    .io_portA_write_data_28(mem_io_portA_write_data_28),
    .io_portA_write_data_29(mem_io_portA_write_data_29),
    .io_portA_write_data_30(mem_io_portA_write_data_30),
    .io_portA_write_data_31(mem_io_portA_write_data_31),
    .io_portB_address(mem_io_portB_address),
    .io_portB_read_enable(mem_io_portB_read_enable),
    .io_portB_read_data_0(mem_io_portB_read_data_0),
    .io_portB_read_data_1(mem_io_portB_read_data_1),
    .io_portB_read_data_2(mem_io_portB_read_data_2),
    .io_portB_read_data_3(mem_io_portB_read_data_3),
    .io_portB_read_data_4(mem_io_portB_read_data_4),
    .io_portB_read_data_5(mem_io_portB_read_data_5),
    .io_portB_read_data_6(mem_io_portB_read_data_6),
    .io_portB_read_data_7(mem_io_portB_read_data_7),
    .io_portB_read_data_8(mem_io_portB_read_data_8),
    .io_portB_read_data_9(mem_io_portB_read_data_9),
    .io_portB_read_data_10(mem_io_portB_read_data_10),
    .io_portB_read_data_11(mem_io_portB_read_data_11),
    .io_portB_read_data_12(mem_io_portB_read_data_12),
    .io_portB_read_data_13(mem_io_portB_read_data_13),
    .io_portB_read_data_14(mem_io_portB_read_data_14),
    .io_portB_read_data_15(mem_io_portB_read_data_15),
    .io_portB_read_data_16(mem_io_portB_read_data_16),
    .io_portB_read_data_17(mem_io_portB_read_data_17),
    .io_portB_read_data_18(mem_io_portB_read_data_18),
    .io_portB_read_data_19(mem_io_portB_read_data_19),
    .io_portB_read_data_20(mem_io_portB_read_data_20),
    .io_portB_read_data_21(mem_io_portB_read_data_21),
    .io_portB_read_data_22(mem_io_portB_read_data_22),
    .io_portB_read_data_23(mem_io_portB_read_data_23),
    .io_portB_read_data_24(mem_io_portB_read_data_24),
    .io_portB_read_data_25(mem_io_portB_read_data_25),
    .io_portB_read_data_26(mem_io_portB_read_data_26),
    .io_portB_read_data_27(mem_io_portB_read_data_27),
    .io_portB_read_data_28(mem_io_portB_read_data_28),
    .io_portB_read_data_29(mem_io_portB_read_data_29),
    .io_portB_read_data_30(mem_io_portB_read_data_30),
    .io_portB_read_data_31(mem_io_portB_read_data_31),
    .io_portB_write_enable(mem_io_portB_write_enable),
    .io_portB_write_data_0(mem_io_portB_write_data_0),
    .io_portB_write_data_1(mem_io_portB_write_data_1),
    .io_portB_write_data_2(mem_io_portB_write_data_2),
    .io_portB_write_data_3(mem_io_portB_write_data_3),
    .io_portB_write_data_4(mem_io_portB_write_data_4),
    .io_portB_write_data_5(mem_io_portB_write_data_5),
    .io_portB_write_data_6(mem_io_portB_write_data_6),
    .io_portB_write_data_7(mem_io_portB_write_data_7),
    .io_portB_write_data_8(mem_io_portB_write_data_8),
    .io_portB_write_data_9(mem_io_portB_write_data_9),
    .io_portB_write_data_10(mem_io_portB_write_data_10),
    .io_portB_write_data_11(mem_io_portB_write_data_11),
    .io_portB_write_data_12(mem_io_portB_write_data_12),
    .io_portB_write_data_13(mem_io_portB_write_data_13),
    .io_portB_write_data_14(mem_io_portB_write_data_14),
    .io_portB_write_data_15(mem_io_portB_write_data_15),
    .io_portB_write_data_16(mem_io_portB_write_data_16),
    .io_portB_write_data_17(mem_io_portB_write_data_17),
    .io_portB_write_data_18(mem_io_portB_write_data_18),
    .io_portB_write_data_19(mem_io_portB_write_data_19),
    .io_portB_write_data_20(mem_io_portB_write_data_20),
    .io_portB_write_data_21(mem_io_portB_write_data_21),
    .io_portB_write_data_22(mem_io_portB_write_data_22),
    .io_portB_write_data_23(mem_io_portB_write_data_23),
    .io_portB_write_data_24(mem_io_portB_write_data_24),
    .io_portB_write_data_25(mem_io_portB_write_data_25),
    .io_portB_write_data_26(mem_io_portB_write_data_26),
    .io_portB_write_data_27(mem_io_portB_write_data_27),
    .io_portB_write_data_28(mem_io_portB_write_data_28),
    .io_portB_write_data_29(mem_io_portB_write_data_29),
    .io_portB_write_data_30(mem_io_portB_write_data_30),
    .io_portB_write_data_31(mem_io_portB_write_data_31)
  );
  Queue_10 output_ ( // @[DualPortMem.scala 48:24]
    .clock(output__clock),
    .reset(output__reset),
    .io_enq_ready(output__io_enq_ready),
    .io_enq_valid(output__io_enq_valid),
    .io_enq_bits_0(output__io_enq_bits_0),
    .io_enq_bits_1(output__io_enq_bits_1),
    .io_enq_bits_2(output__io_enq_bits_2),
    .io_enq_bits_3(output__io_enq_bits_3),
    .io_enq_bits_4(output__io_enq_bits_4),
    .io_enq_bits_5(output__io_enq_bits_5),
    .io_enq_bits_6(output__io_enq_bits_6),
    .io_enq_bits_7(output__io_enq_bits_7),
    .io_enq_bits_8(output__io_enq_bits_8),
    .io_enq_bits_9(output__io_enq_bits_9),
    .io_enq_bits_10(output__io_enq_bits_10),
    .io_enq_bits_11(output__io_enq_bits_11),
    .io_enq_bits_12(output__io_enq_bits_12),
    .io_enq_bits_13(output__io_enq_bits_13),
    .io_enq_bits_14(output__io_enq_bits_14),
    .io_enq_bits_15(output__io_enq_bits_15),
    .io_enq_bits_16(output__io_enq_bits_16),
    .io_enq_bits_17(output__io_enq_bits_17),
    .io_enq_bits_18(output__io_enq_bits_18),
    .io_enq_bits_19(output__io_enq_bits_19),
    .io_enq_bits_20(output__io_enq_bits_20),
    .io_enq_bits_21(output__io_enq_bits_21),
    .io_enq_bits_22(output__io_enq_bits_22),
    .io_enq_bits_23(output__io_enq_bits_23),
    .io_enq_bits_24(output__io_enq_bits_24),
    .io_enq_bits_25(output__io_enq_bits_25),
    .io_enq_bits_26(output__io_enq_bits_26),
    .io_enq_bits_27(output__io_enq_bits_27),
    .io_enq_bits_28(output__io_enq_bits_28),
    .io_enq_bits_29(output__io_enq_bits_29),
    .io_enq_bits_30(output__io_enq_bits_30),
    .io_enq_bits_31(output__io_enq_bits_31),
    .io_deq_ready(output__io_deq_ready),
    .io_deq_valid(output__io_deq_valid),
    .io_deq_bits_0(output__io_deq_bits_0),
    .io_deq_bits_1(output__io_deq_bits_1),
    .io_deq_bits_2(output__io_deq_bits_2),
    .io_deq_bits_3(output__io_deq_bits_3),
    .io_deq_bits_4(output__io_deq_bits_4),
    .io_deq_bits_5(output__io_deq_bits_5),
    .io_deq_bits_6(output__io_deq_bits_6),
    .io_deq_bits_7(output__io_deq_bits_7),
    .io_deq_bits_8(output__io_deq_bits_8),
    .io_deq_bits_9(output__io_deq_bits_9),
    .io_deq_bits_10(output__io_deq_bits_10),
    .io_deq_bits_11(output__io_deq_bits_11),
    .io_deq_bits_12(output__io_deq_bits_12),
    .io_deq_bits_13(output__io_deq_bits_13),
    .io_deq_bits_14(output__io_deq_bits_14),
    .io_deq_bits_15(output__io_deq_bits_15),
    .io_deq_bits_16(output__io_deq_bits_16),
    .io_deq_bits_17(output__io_deq_bits_17),
    .io_deq_bits_18(output__io_deq_bits_18),
    .io_deq_bits_19(output__io_deq_bits_19),
    .io_deq_bits_20(output__io_deq_bits_20),
    .io_deq_bits_21(output__io_deq_bits_21),
    .io_deq_bits_22(output__io_deq_bits_22),
    .io_deq_bits_23(output__io_deq_bits_23),
    .io_deq_bits_24(output__io_deq_bits_24),
    .io_deq_bits_25(output__io_deq_bits_25),
    .io_deq_bits_26(output__io_deq_bits_26),
    .io_deq_bits_27(output__io_deq_bits_27),
    .io_deq_bits_28(output__io_deq_bits_28),
    .io_deq_bits_29(output__io_deq_bits_29),
    .io_deq_bits_30(output__io_deq_bits_30),
    .io_deq_bits_31(output__io_deq_bits_31),
    .io_count(output__io_count)
  );
  Queue_10 output_1 ( // @[DualPortMem.scala 48:24]
    .clock(output_1_clock),
    .reset(output_1_reset),
    .io_enq_ready(output_1_io_enq_ready),
    .io_enq_valid(output_1_io_enq_valid),
    .io_enq_bits_0(output_1_io_enq_bits_0),
    .io_enq_bits_1(output_1_io_enq_bits_1),
    .io_enq_bits_2(output_1_io_enq_bits_2),
    .io_enq_bits_3(output_1_io_enq_bits_3),
    .io_enq_bits_4(output_1_io_enq_bits_4),
    .io_enq_bits_5(output_1_io_enq_bits_5),
    .io_enq_bits_6(output_1_io_enq_bits_6),
    .io_enq_bits_7(output_1_io_enq_bits_7),
    .io_enq_bits_8(output_1_io_enq_bits_8),
    .io_enq_bits_9(output_1_io_enq_bits_9),
    .io_enq_bits_10(output_1_io_enq_bits_10),
    .io_enq_bits_11(output_1_io_enq_bits_11),
    .io_enq_bits_12(output_1_io_enq_bits_12),
    .io_enq_bits_13(output_1_io_enq_bits_13),
    .io_enq_bits_14(output_1_io_enq_bits_14),
    .io_enq_bits_15(output_1_io_enq_bits_15),
    .io_enq_bits_16(output_1_io_enq_bits_16),
    .io_enq_bits_17(output_1_io_enq_bits_17),
    .io_enq_bits_18(output_1_io_enq_bits_18),
    .io_enq_bits_19(output_1_io_enq_bits_19),
    .io_enq_bits_20(output_1_io_enq_bits_20),
    .io_enq_bits_21(output_1_io_enq_bits_21),
    .io_enq_bits_22(output_1_io_enq_bits_22),
    .io_enq_bits_23(output_1_io_enq_bits_23),
    .io_enq_bits_24(output_1_io_enq_bits_24),
    .io_enq_bits_25(output_1_io_enq_bits_25),
    .io_enq_bits_26(output_1_io_enq_bits_26),
    .io_enq_bits_27(output_1_io_enq_bits_27),
    .io_enq_bits_28(output_1_io_enq_bits_28),
    .io_enq_bits_29(output_1_io_enq_bits_29),
    .io_enq_bits_30(output_1_io_enq_bits_30),
    .io_enq_bits_31(output_1_io_enq_bits_31),
    .io_deq_ready(output_1_io_deq_ready),
    .io_deq_valid(output_1_io_deq_valid),
    .io_deq_bits_0(output_1_io_deq_bits_0),
    .io_deq_bits_1(output_1_io_deq_bits_1),
    .io_deq_bits_2(output_1_io_deq_bits_2),
    .io_deq_bits_3(output_1_io_deq_bits_3),
    .io_deq_bits_4(output_1_io_deq_bits_4),
    .io_deq_bits_5(output_1_io_deq_bits_5),
    .io_deq_bits_6(output_1_io_deq_bits_6),
    .io_deq_bits_7(output_1_io_deq_bits_7),
    .io_deq_bits_8(output_1_io_deq_bits_8),
    .io_deq_bits_9(output_1_io_deq_bits_9),
    .io_deq_bits_10(output_1_io_deq_bits_10),
    .io_deq_bits_11(output_1_io_deq_bits_11),
    .io_deq_bits_12(output_1_io_deq_bits_12),
    .io_deq_bits_13(output_1_io_deq_bits_13),
    .io_deq_bits_14(output_1_io_deq_bits_14),
    .io_deq_bits_15(output_1_io_deq_bits_15),
    .io_deq_bits_16(output_1_io_deq_bits_16),
    .io_deq_bits_17(output_1_io_deq_bits_17),
    .io_deq_bits_18(output_1_io_deq_bits_18),
    .io_deq_bits_19(output_1_io_deq_bits_19),
    .io_deq_bits_20(output_1_io_deq_bits_20),
    .io_deq_bits_21(output_1_io_deq_bits_21),
    .io_deq_bits_22(output_1_io_deq_bits_22),
    .io_deq_bits_23(output_1_io_deq_bits_23),
    .io_deq_bits_24(output_1_io_deq_bits_24),
    .io_deq_bits_25(output_1_io_deq_bits_25),
    .io_deq_bits_26(output_1_io_deq_bits_26),
    .io_deq_bits_27(output_1_io_deq_bits_27),
    .io_deq_bits_28(output_1_io_deq_bits_28),
    .io_deq_bits_29(output_1_io_deq_bits_29),
    .io_deq_bits_30(output_1_io_deq_bits_30),
    .io_deq_bits_31(output_1_io_deq_bits_31),
    .io_count(output_1_io_count)
  );
  assign io_portA_control_ready = io_portA_control_bits_write ? io_portA_input_valid : outputReady; // @[DualPortMem.scala 59:30 60:21 64:21]
  assign io_portA_input_ready = io_portA_control_valid & io_portA_control_bits_write; // @[DualPortMem.scala 75:34]
  assign io_portA_output_valid = output__io_deq_valid; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_0 = output__io_deq_bits_0; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_1 = output__io_deq_bits_1; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_2 = output__io_deq_bits_2; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_3 = output__io_deq_bits_3; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_4 = output__io_deq_bits_4; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_5 = output__io_deq_bits_5; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_6 = output__io_deq_bits_6; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_7 = output__io_deq_bits_7; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_8 = output__io_deq_bits_8; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_9 = output__io_deq_bits_9; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_10 = output__io_deq_bits_10; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_11 = output__io_deq_bits_11; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_12 = output__io_deq_bits_12; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_13 = output__io_deq_bits_13; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_14 = output__io_deq_bits_14; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_15 = output__io_deq_bits_15; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_16 = output__io_deq_bits_16; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_17 = output__io_deq_bits_17; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_18 = output__io_deq_bits_18; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_19 = output__io_deq_bits_19; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_20 = output__io_deq_bits_20; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_21 = output__io_deq_bits_21; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_22 = output__io_deq_bits_22; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_23 = output__io_deq_bits_23; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_24 = output__io_deq_bits_24; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_25 = output__io_deq_bits_25; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_26 = output__io_deq_bits_26; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_27 = output__io_deq_bits_27; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_28 = output__io_deq_bits_28; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_29 = output__io_deq_bits_29; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_30 = output__io_deq_bits_30; // @[DualPortMem.scala 72:17]
  assign io_portA_output_bits_31 = output__io_deq_bits_31; // @[DualPortMem.scala 72:17]
  assign io_portB_control_ready = io_portB_control_bits_write ? io_portB_input_valid : outputReady_1; // @[DualPortMem.scala 59:30 60:21 64:21]
  assign io_portB_input_ready = io_portB_control_valid & io_portB_control_bits_write; // @[DualPortMem.scala 75:34]
  assign io_portB_output_valid = output_1_io_deq_valid; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_0 = output_1_io_deq_bits_0; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_1 = output_1_io_deq_bits_1; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_2 = output_1_io_deq_bits_2; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_3 = output_1_io_deq_bits_3; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_4 = output_1_io_deq_bits_4; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_5 = output_1_io_deq_bits_5; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_6 = output_1_io_deq_bits_6; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_7 = output_1_io_deq_bits_7; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_8 = output_1_io_deq_bits_8; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_9 = output_1_io_deq_bits_9; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_10 = output_1_io_deq_bits_10; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_11 = output_1_io_deq_bits_11; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_12 = output_1_io_deq_bits_12; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_13 = output_1_io_deq_bits_13; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_14 = output_1_io_deq_bits_14; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_15 = output_1_io_deq_bits_15; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_16 = output_1_io_deq_bits_16; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_17 = output_1_io_deq_bits_17; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_18 = output_1_io_deq_bits_18; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_19 = output_1_io_deq_bits_19; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_20 = output_1_io_deq_bits_20; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_21 = output_1_io_deq_bits_21; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_22 = output_1_io_deq_bits_22; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_23 = output_1_io_deq_bits_23; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_24 = output_1_io_deq_bits_24; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_25 = output_1_io_deq_bits_25; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_26 = output_1_io_deq_bits_26; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_27 = output_1_io_deq_bits_27; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_28 = output_1_io_deq_bits_28; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_29 = output_1_io_deq_bits_29; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_30 = output_1_io_deq_bits_30; // @[DualPortMem.scala 72:17]
  assign io_portB_output_bits_31 = output_1_io_deq_bits_31; // @[DualPortMem.scala 72:17]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_portA_address = io_portA_control_bits_address; // @[DualPortMem.scala 57:19]
  assign mem_io_portA_read_enable = io_portA_control_bits_write ? 1'h0 : io_portA_control_valid & outputReady; // @[DualPortMem.scala 59:30 62:25 66:25]
  assign mem_io_portA_write_enable = io_portA_control_bits_write & (io_portA_control_valid & io_portA_input_valid); // @[DualPortMem.scala 59:30 61:26 65:26]
  assign mem_io_portA_write_data_0 = io_portA_input_bits_0; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_1 = io_portA_input_bits_1; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_2 = io_portA_input_bits_2; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_3 = io_portA_input_bits_3; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_4 = io_portA_input_bits_4; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_5 = io_portA_input_bits_5; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_6 = io_portA_input_bits_6; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_7 = io_portA_input_bits_7; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_8 = io_portA_input_bits_8; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_9 = io_portA_input_bits_9; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_10 = io_portA_input_bits_10; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_11 = io_portA_input_bits_11; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_12 = io_portA_input_bits_12; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_13 = io_portA_input_bits_13; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_14 = io_portA_input_bits_14; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_15 = io_portA_input_bits_15; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_16 = io_portA_input_bits_16; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_17 = io_portA_input_bits_17; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_18 = io_portA_input_bits_18; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_19 = io_portA_input_bits_19; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_20 = io_portA_input_bits_20; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_21 = io_portA_input_bits_21; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_22 = io_portA_input_bits_22; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_23 = io_portA_input_bits_23; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_24 = io_portA_input_bits_24; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_25 = io_portA_input_bits_25; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_26 = io_portA_input_bits_26; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_27 = io_portA_input_bits_27; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_28 = io_portA_input_bits_28; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_29 = io_portA_input_bits_29; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_30 = io_portA_input_bits_30; // @[DualPortMem.scala 74:22]
  assign mem_io_portA_write_data_31 = io_portA_input_bits_31; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_address = io_portB_control_bits_address; // @[DualPortMem.scala 57:19]
  assign mem_io_portB_read_enable = io_portB_control_bits_write ? 1'h0 : io_portB_control_valid & outputReady_1; // @[DualPortMem.scala 59:30 62:25 66:25]
  assign mem_io_portB_write_enable = io_portB_control_bits_write & (io_portB_control_valid & io_portB_input_valid); // @[DualPortMem.scala 59:30 61:26 65:26]
  assign mem_io_portB_write_data_0 = io_portB_input_bits_0; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_1 = io_portB_input_bits_1; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_2 = io_portB_input_bits_2; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_3 = io_portB_input_bits_3; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_4 = io_portB_input_bits_4; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_5 = io_portB_input_bits_5; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_6 = io_portB_input_bits_6; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_7 = io_portB_input_bits_7; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_8 = io_portB_input_bits_8; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_9 = io_portB_input_bits_9; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_10 = io_portB_input_bits_10; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_11 = io_portB_input_bits_11; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_12 = io_portB_input_bits_12; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_13 = io_portB_input_bits_13; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_14 = io_portB_input_bits_14; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_15 = io_portB_input_bits_15; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_16 = io_portB_input_bits_16; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_17 = io_portB_input_bits_17; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_18 = io_portB_input_bits_18; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_19 = io_portB_input_bits_19; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_20 = io_portB_input_bits_20; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_21 = io_portB_input_bits_21; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_22 = io_portB_input_bits_22; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_23 = io_portB_input_bits_23; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_24 = io_portB_input_bits_24; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_25 = io_portB_input_bits_25; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_26 = io_portB_input_bits_26; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_27 = io_portB_input_bits_27; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_28 = io_portB_input_bits_28; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_29 = io_portB_input_bits_29; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_30 = io_portB_input_bits_30; // @[DualPortMem.scala 74:22]
  assign mem_io_portB_write_data_31 = io_portB_input_bits_31; // @[DualPortMem.scala 74:22]
  assign output__clock = clock;
  assign output__reset = reset;
  assign output__io_enq_valid = output_io_enq_valid_sr_0; // @[DualPortMem.scala 70:25]
  assign output__io_enq_bits_0 = mem_io_portA_read_data_0; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_1 = mem_io_portA_read_data_1; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_2 = mem_io_portA_read_data_2; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_3 = mem_io_portA_read_data_3; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_4 = mem_io_portA_read_data_4; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_5 = mem_io_portA_read_data_5; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_6 = mem_io_portA_read_data_6; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_7 = mem_io_portA_read_data_7; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_8 = mem_io_portA_read_data_8; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_9 = mem_io_portA_read_data_9; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_10 = mem_io_portA_read_data_10; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_11 = mem_io_portA_read_data_11; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_12 = mem_io_portA_read_data_12; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_13 = mem_io_portA_read_data_13; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_14 = mem_io_portA_read_data_14; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_15 = mem_io_portA_read_data_15; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_16 = mem_io_portA_read_data_16; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_17 = mem_io_portA_read_data_17; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_18 = mem_io_portA_read_data_18; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_19 = mem_io_portA_read_data_19; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_20 = mem_io_portA_read_data_20; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_21 = mem_io_portA_read_data_21; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_22 = mem_io_portA_read_data_22; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_23 = mem_io_portA_read_data_23; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_24 = mem_io_portA_read_data_24; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_25 = mem_io_portA_read_data_25; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_26 = mem_io_portA_read_data_26; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_27 = mem_io_portA_read_data_27; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_28 = mem_io_portA_read_data_28; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_29 = mem_io_portA_read_data_29; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_30 = mem_io_portA_read_data_30; // @[DualPortMem.scala 69:24]
  assign output__io_enq_bits_31 = mem_io_portA_read_data_31; // @[DualPortMem.scala 69:24]
  assign output__io_deq_ready = io_portA_output_ready; // @[DualPortMem.scala 72:17]
  assign output_1_clock = clock;
  assign output_1_reset = reset;
  assign output_1_io_enq_valid = output_io_enq_valid_sr_1_0; // @[DualPortMem.scala 70:25]
  assign output_1_io_enq_bits_0 = mem_io_portB_read_data_0; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_1 = mem_io_portB_read_data_1; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_2 = mem_io_portB_read_data_2; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_3 = mem_io_portB_read_data_3; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_4 = mem_io_portB_read_data_4; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_5 = mem_io_portB_read_data_5; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_6 = mem_io_portB_read_data_6; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_7 = mem_io_portB_read_data_7; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_8 = mem_io_portB_read_data_8; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_9 = mem_io_portB_read_data_9; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_10 = mem_io_portB_read_data_10; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_11 = mem_io_portB_read_data_11; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_12 = mem_io_portB_read_data_12; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_13 = mem_io_portB_read_data_13; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_14 = mem_io_portB_read_data_14; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_15 = mem_io_portB_read_data_15; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_16 = mem_io_portB_read_data_16; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_17 = mem_io_portB_read_data_17; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_18 = mem_io_portB_read_data_18; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_19 = mem_io_portB_read_data_19; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_20 = mem_io_portB_read_data_20; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_21 = mem_io_portB_read_data_21; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_22 = mem_io_portB_read_data_22; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_23 = mem_io_portB_read_data_23; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_24 = mem_io_portB_read_data_24; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_25 = mem_io_portB_read_data_25; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_26 = mem_io_portB_read_data_26; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_27 = mem_io_portB_read_data_27; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_28 = mem_io_portB_read_data_28; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_29 = mem_io_portB_read_data_29; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_30 = mem_io_portB_read_data_30; // @[DualPortMem.scala 69:24]
  assign output_1_io_enq_bits_31 = mem_io_portB_read_data_31; // @[DualPortMem.scala 69:24]
  assign output_1_io_deq_ready = io_portB_output_ready; // @[DualPortMem.scala 72:17]
  always @(posedge clock) begin
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_0 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_0 <= mem_io_portA_read_enable; // @[ShiftRegister.scala 25:12]
    end
    if (reset) begin // @[ShiftRegister.scala 10:22]
      output_io_enq_valid_sr_1_0 <= 1'h0; // @[ShiftRegister.scala 10:22]
    end else begin
      output_io_enq_valid_sr_1_0 <= mem_io_portB_read_enable; // @[ShiftRegister.scala 25:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  output_io_enq_valid_sr_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  output_io_enq_valid_sr_1_0 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Demux_3(
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_0,
  input  [15:0] io_in_bits_1,
  input  [15:0] io_in_bits_2,
  input  [15:0] io_in_bits_3,
  input  [15:0] io_in_bits_4,
  input  [15:0] io_in_bits_5,
  input  [15:0] io_in_bits_6,
  input  [15:0] io_in_bits_7,
  input  [15:0] io_in_bits_8,
  input  [15:0] io_in_bits_9,
  input  [15:0] io_in_bits_10,
  input  [15:0] io_in_bits_11,
  input  [15:0] io_in_bits_12,
  input  [15:0] io_in_bits_13,
  input  [15:0] io_in_bits_14,
  input  [15:0] io_in_bits_15,
  input  [15:0] io_in_bits_16,
  input  [15:0] io_in_bits_17,
  input  [15:0] io_in_bits_18,
  input  [15:0] io_in_bits_19,
  input  [15:0] io_in_bits_20,
  input  [15:0] io_in_bits_21,
  input  [15:0] io_in_bits_22,
  input  [15:0] io_in_bits_23,
  input  [15:0] io_in_bits_24,
  input  [15:0] io_in_bits_25,
  input  [15:0] io_in_bits_26,
  input  [15:0] io_in_bits_27,
  input  [15:0] io_in_bits_28,
  input  [15:0] io_in_bits_29,
  input  [15:0] io_in_bits_30,
  input  [15:0] io_in_bits_31,
  output        io_sel_ready,
  input         io_sel_valid,
  input  [1:0]  io_sel_bits,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [15:0] io_out_0_bits_0,
  output [15:0] io_out_0_bits_1,
  output [15:0] io_out_0_bits_2,
  output [15:0] io_out_0_bits_3,
  output [15:0] io_out_0_bits_4,
  output [15:0] io_out_0_bits_5,
  output [15:0] io_out_0_bits_6,
  output [15:0] io_out_0_bits_7,
  output [15:0] io_out_0_bits_8,
  output [15:0] io_out_0_bits_9,
  output [15:0] io_out_0_bits_10,
  output [15:0] io_out_0_bits_11,
  output [15:0] io_out_0_bits_12,
  output [15:0] io_out_0_bits_13,
  output [15:0] io_out_0_bits_14,
  output [15:0] io_out_0_bits_15,
  output [15:0] io_out_0_bits_16,
  output [15:0] io_out_0_bits_17,
  output [15:0] io_out_0_bits_18,
  output [15:0] io_out_0_bits_19,
  output [15:0] io_out_0_bits_20,
  output [15:0] io_out_0_bits_21,
  output [15:0] io_out_0_bits_22,
  output [15:0] io_out_0_bits_23,
  output [15:0] io_out_0_bits_24,
  output [15:0] io_out_0_bits_25,
  output [15:0] io_out_0_bits_26,
  output [15:0] io_out_0_bits_27,
  output [15:0] io_out_0_bits_28,
  output [15:0] io_out_0_bits_29,
  output [15:0] io_out_0_bits_30,
  output [15:0] io_out_0_bits_31,
  input         io_out_1_ready,
  output        io_out_1_valid,
  output [15:0] io_out_1_bits_0,
  output [15:0] io_out_1_bits_1,
  output [15:0] io_out_1_bits_2,
  output [15:0] io_out_1_bits_3,
  output [15:0] io_out_1_bits_4,
  output [15:0] io_out_1_bits_5,
  output [15:0] io_out_1_bits_6,
  output [15:0] io_out_1_bits_7,
  output [15:0] io_out_1_bits_8,
  output [15:0] io_out_1_bits_9,
  output [15:0] io_out_1_bits_10,
  output [15:0] io_out_1_bits_11,
  output [15:0] io_out_1_bits_12,
  output [15:0] io_out_1_bits_13,
  output [15:0] io_out_1_bits_14,
  output [15:0] io_out_1_bits_15,
  output [15:0] io_out_1_bits_16,
  output [15:0] io_out_1_bits_17,
  output [15:0] io_out_1_bits_18,
  output [15:0] io_out_1_bits_19,
  output [15:0] io_out_1_bits_20,
  output [15:0] io_out_1_bits_21,
  output [15:0] io_out_1_bits_22,
  output [15:0] io_out_1_bits_23,
  output [15:0] io_out_1_bits_24,
  output [15:0] io_out_1_bits_25,
  output [15:0] io_out_1_bits_26,
  output [15:0] io_out_1_bits_27,
  output [15:0] io_out_1_bits_28,
  output [15:0] io_out_1_bits_29,
  output [15:0] io_out_1_bits_30,
  output [15:0] io_out_1_bits_31,
  input         io_out_2_ready,
  output        io_out_2_valid,
  output [15:0] io_out_2_bits_0,
  output [15:0] io_out_2_bits_1,
  output [15:0] io_out_2_bits_2,
  output [15:0] io_out_2_bits_3,
  output [15:0] io_out_2_bits_4,
  output [15:0] io_out_2_bits_5,
  output [15:0] io_out_2_bits_6,
  output [15:0] io_out_2_bits_7,
  output [15:0] io_out_2_bits_8,
  output [15:0] io_out_2_bits_9,
  output [15:0] io_out_2_bits_10,
  output [15:0] io_out_2_bits_11,
  output [15:0] io_out_2_bits_12,
  output [15:0] io_out_2_bits_13,
  output [15:0] io_out_2_bits_14,
  output [15:0] io_out_2_bits_15,
  output [15:0] io_out_2_bits_16,
  output [15:0] io_out_2_bits_17,
  output [15:0] io_out_2_bits_18,
  output [15:0] io_out_2_bits_19,
  output [15:0] io_out_2_bits_20,
  output [15:0] io_out_2_bits_21,
  output [15:0] io_out_2_bits_22,
  output [15:0] io_out_2_bits_23,
  output [15:0] io_out_2_bits_24,
  output [15:0] io_out_2_bits_25,
  output [15:0] io_out_2_bits_26,
  output [15:0] io_out_2_bits_27,
  output [15:0] io_out_2_bits_28,
  output [15:0] io_out_2_bits_29,
  output [15:0] io_out_2_bits_30,
  output [15:0] io_out_2_bits_31
);
  wire  _GEN_100 = 2'h1 == io_sel_bits ? io_out_1_ready : io_out_0_ready; // @[Demux.scala 34:{25,25}]
  wire  _GEN_101 = 2'h2 == io_sel_bits ? io_out_2_ready : _GEN_100; // @[Demux.scala 34:{25,25}]
  assign io_in_ready = io_sel_valid & _GEN_101; // @[Demux.scala 35:25]
  assign io_sel_ready = io_in_valid & _GEN_101; // @[Demux.scala 34:25]
  assign io_out_0_valid = 2'h0 == io_sel_bits & (io_sel_valid & io_in_valid); // @[Demux.scala 33:{13,13} 28:15]
  assign io_out_0_bits_0 = 2'h0 == io_sel_bits ? $signed(io_in_bits_0) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_1 = 2'h0 == io_sel_bits ? $signed(io_in_bits_1) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_2 = 2'h0 == io_sel_bits ? $signed(io_in_bits_2) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_3 = 2'h0 == io_sel_bits ? $signed(io_in_bits_3) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_4 = 2'h0 == io_sel_bits ? $signed(io_in_bits_4) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_5 = 2'h0 == io_sel_bits ? $signed(io_in_bits_5) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_6 = 2'h0 == io_sel_bits ? $signed(io_in_bits_6) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_7 = 2'h0 == io_sel_bits ? $signed(io_in_bits_7) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_8 = 2'h0 == io_sel_bits ? $signed(io_in_bits_8) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_9 = 2'h0 == io_sel_bits ? $signed(io_in_bits_9) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_10 = 2'h0 == io_sel_bits ? $signed(io_in_bits_10) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_11 = 2'h0 == io_sel_bits ? $signed(io_in_bits_11) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_12 = 2'h0 == io_sel_bits ? $signed(io_in_bits_12) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_13 = 2'h0 == io_sel_bits ? $signed(io_in_bits_13) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_14 = 2'h0 == io_sel_bits ? $signed(io_in_bits_14) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_15 = 2'h0 == io_sel_bits ? $signed(io_in_bits_15) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_16 = 2'h0 == io_sel_bits ? $signed(io_in_bits_16) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_17 = 2'h0 == io_sel_bits ? $signed(io_in_bits_17) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_18 = 2'h0 == io_sel_bits ? $signed(io_in_bits_18) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_19 = 2'h0 == io_sel_bits ? $signed(io_in_bits_19) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_20 = 2'h0 == io_sel_bits ? $signed(io_in_bits_20) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_21 = 2'h0 == io_sel_bits ? $signed(io_in_bits_21) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_22 = 2'h0 == io_sel_bits ? $signed(io_in_bits_22) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_23 = 2'h0 == io_sel_bits ? $signed(io_in_bits_23) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_24 = 2'h0 == io_sel_bits ? $signed(io_in_bits_24) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_25 = 2'h0 == io_sel_bits ? $signed(io_in_bits_25) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_26 = 2'h0 == io_sel_bits ? $signed(io_in_bits_26) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_27 = 2'h0 == io_sel_bits ? $signed(io_in_bits_27) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_28 = 2'h0 == io_sel_bits ? $signed(io_in_bits_28) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_29 = 2'h0 == io_sel_bits ? $signed(io_in_bits_29) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_30 = 2'h0 == io_sel_bits ? $signed(io_in_bits_30) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_0_bits_31 = 2'h0 == io_sel_bits ? $signed(io_in_bits_31) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_valid = 2'h1 == io_sel_bits & (io_sel_valid & io_in_valid); // @[Demux.scala 33:{13,13} 28:15]
  assign io_out_1_bits_0 = 2'h1 == io_sel_bits ? $signed(io_in_bits_0) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_1 = 2'h1 == io_sel_bits ? $signed(io_in_bits_1) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_2 = 2'h1 == io_sel_bits ? $signed(io_in_bits_2) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_3 = 2'h1 == io_sel_bits ? $signed(io_in_bits_3) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_4 = 2'h1 == io_sel_bits ? $signed(io_in_bits_4) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_5 = 2'h1 == io_sel_bits ? $signed(io_in_bits_5) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_6 = 2'h1 == io_sel_bits ? $signed(io_in_bits_6) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_7 = 2'h1 == io_sel_bits ? $signed(io_in_bits_7) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_8 = 2'h1 == io_sel_bits ? $signed(io_in_bits_8) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_9 = 2'h1 == io_sel_bits ? $signed(io_in_bits_9) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_10 = 2'h1 == io_sel_bits ? $signed(io_in_bits_10) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_11 = 2'h1 == io_sel_bits ? $signed(io_in_bits_11) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_12 = 2'h1 == io_sel_bits ? $signed(io_in_bits_12) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_13 = 2'h1 == io_sel_bits ? $signed(io_in_bits_13) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_14 = 2'h1 == io_sel_bits ? $signed(io_in_bits_14) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_15 = 2'h1 == io_sel_bits ? $signed(io_in_bits_15) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_16 = 2'h1 == io_sel_bits ? $signed(io_in_bits_16) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_17 = 2'h1 == io_sel_bits ? $signed(io_in_bits_17) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_18 = 2'h1 == io_sel_bits ? $signed(io_in_bits_18) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_19 = 2'h1 == io_sel_bits ? $signed(io_in_bits_19) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_20 = 2'h1 == io_sel_bits ? $signed(io_in_bits_20) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_21 = 2'h1 == io_sel_bits ? $signed(io_in_bits_21) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_22 = 2'h1 == io_sel_bits ? $signed(io_in_bits_22) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_23 = 2'h1 == io_sel_bits ? $signed(io_in_bits_23) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_24 = 2'h1 == io_sel_bits ? $signed(io_in_bits_24) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_25 = 2'h1 == io_sel_bits ? $signed(io_in_bits_25) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_26 = 2'h1 == io_sel_bits ? $signed(io_in_bits_26) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_27 = 2'h1 == io_sel_bits ? $signed(io_in_bits_27) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_28 = 2'h1 == io_sel_bits ? $signed(io_in_bits_28) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_29 = 2'h1 == io_sel_bits ? $signed(io_in_bits_29) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_30 = 2'h1 == io_sel_bits ? $signed(io_in_bits_30) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_1_bits_31 = 2'h1 == io_sel_bits ? $signed(io_in_bits_31) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_valid = 2'h2 == io_sel_bits & (io_sel_valid & io_in_valid); // @[Demux.scala 33:{13,13} 28:15]
  assign io_out_2_bits_0 = 2'h2 == io_sel_bits ? $signed(io_in_bits_0) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_1 = 2'h2 == io_sel_bits ? $signed(io_in_bits_1) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_2 = 2'h2 == io_sel_bits ? $signed(io_in_bits_2) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_3 = 2'h2 == io_sel_bits ? $signed(io_in_bits_3) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_4 = 2'h2 == io_sel_bits ? $signed(io_in_bits_4) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_5 = 2'h2 == io_sel_bits ? $signed(io_in_bits_5) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_6 = 2'h2 == io_sel_bits ? $signed(io_in_bits_6) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_7 = 2'h2 == io_sel_bits ? $signed(io_in_bits_7) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_8 = 2'h2 == io_sel_bits ? $signed(io_in_bits_8) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_9 = 2'h2 == io_sel_bits ? $signed(io_in_bits_9) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_10 = 2'h2 == io_sel_bits ? $signed(io_in_bits_10) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_11 = 2'h2 == io_sel_bits ? $signed(io_in_bits_11) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_12 = 2'h2 == io_sel_bits ? $signed(io_in_bits_12) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_13 = 2'h2 == io_sel_bits ? $signed(io_in_bits_13) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_14 = 2'h2 == io_sel_bits ? $signed(io_in_bits_14) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_15 = 2'h2 == io_sel_bits ? $signed(io_in_bits_15) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_16 = 2'h2 == io_sel_bits ? $signed(io_in_bits_16) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_17 = 2'h2 == io_sel_bits ? $signed(io_in_bits_17) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_18 = 2'h2 == io_sel_bits ? $signed(io_in_bits_18) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_19 = 2'h2 == io_sel_bits ? $signed(io_in_bits_19) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_20 = 2'h2 == io_sel_bits ? $signed(io_in_bits_20) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_21 = 2'h2 == io_sel_bits ? $signed(io_in_bits_21) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_22 = 2'h2 == io_sel_bits ? $signed(io_in_bits_22) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_23 = 2'h2 == io_sel_bits ? $signed(io_in_bits_23) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_24 = 2'h2 == io_sel_bits ? $signed(io_in_bits_24) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_25 = 2'h2 == io_sel_bits ? $signed(io_in_bits_25) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_26 = 2'h2 == io_sel_bits ? $signed(io_in_bits_26) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_27 = 2'h2 == io_sel_bits ? $signed(io_in_bits_27) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_28 = 2'h2 == io_sel_bits ? $signed(io_in_bits_28) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_29 = 2'h2 == io_sel_bits ? $signed(io_in_bits_29) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_30 = 2'h2 == io_sel_bits ? $signed(io_in_bits_30) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
  assign io_out_2_bits_31 = 2'h2 == io_sel_bits ? $signed(io_in_bits_31) : $signed(16'sh0); // @[Demux.scala 32:{12,12} 27:14]
endmodule
module SizeHandler_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [1:0]  io_in_bits_sel,
  input  [13:0] io_in_bits_size,
  input         io_out_ready,
  output        io_out_valid,
  output [1:0]  io_out_bits_sel
);
  wire  sizeCounter_clock; // @[Counter.scala 34:19]
  wire  sizeCounter_reset; // @[Counter.scala 34:19]
  wire  sizeCounter_io_value_ready; // @[Counter.scala 34:19]
  wire [13:0] sizeCounter_io_value_bits; // @[Counter.scala 34:19]
  wire  sizeCounter_io_resetValue; // @[Counter.scala 34:19]
  wire  fire = io_in_valid & io_out_ready; // @[SizeHandler.scala 32:23]
  Counter_2 sizeCounter ( // @[Counter.scala 34:19]
    .clock(sizeCounter_clock),
    .reset(sizeCounter_reset),
    .io_value_ready(sizeCounter_io_value_ready),
    .io_value_bits(sizeCounter_io_value_bits),
    .io_resetValue(sizeCounter_io_resetValue)
  );
  assign io_in_ready = sizeCounter_io_value_bits == io_in_bits_size & io_out_ready; // @[SizeHandler.scala 34:52 35:14 38:14]
  assign io_out_valid = io_in_valid; // @[SizeHandler.scala 25:16]
  assign io_out_bits_sel = io_in_bits_sel; // @[SizeHandler.scala 28:34]
  assign sizeCounter_clock = clock;
  assign sizeCounter_reset = reset;
  assign sizeCounter_io_value_ready = sizeCounter_io_value_bits == io_in_bits_size ? 1'h0 : fire; // @[SizeHandler.scala 34:52 Counter.scala 36:22 SizeHandler.scala 39:32]
  assign sizeCounter_io_resetValue = sizeCounter_io_value_bits == io_in_bits_size & fire; // @[SizeHandler.scala 34:52 Counter.scala 35:21 SizeHandler.scala 36:31]
endmodule
module Queue_25(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_sel,
  input  [13:0] io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_sel,
  output [13:0] io_deq_bits_size
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_sel [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_sel_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_sel_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_sel_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_sel_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_sel_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_sel_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_sel_MPORT_en; // @[Decoupled.scala 259:95]
  reg [13:0] ram_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_10 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_10 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_sel_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sel_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_sel_io_deq_bits_MPORT_data = ram_sel[ram_sel_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_sel_MPORT_data = io_enq_bits_sel;
  assign ram_sel_MPORT_addr = 1'h0;
  assign ram_sel_MPORT_mask = 1'h1;
  assign ram_sel_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_sel = empty ? io_enq_bits_sel : ram_sel_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_sel_MPORT_en & ram_sel_MPORT_mask) begin
      ram_sel[ram_sel_MPORT_addr] <= ram_sel_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_sel[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[13:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SizeHandler_3(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_sel,
  input  [13:0] io_in_bits_size,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_sel
);
  wire  sizeCounter_clock; // @[Counter.scala 34:19]
  wire  sizeCounter_reset; // @[Counter.scala 34:19]
  wire  sizeCounter_io_value_ready; // @[Counter.scala 34:19]
  wire [13:0] sizeCounter_io_value_bits; // @[Counter.scala 34:19]
  wire  sizeCounter_io_resetValue; // @[Counter.scala 34:19]
  wire  fire = io_in_valid & io_out_ready; // @[SizeHandler.scala 32:23]
  Counter_2 sizeCounter ( // @[Counter.scala 34:19]
    .clock(sizeCounter_clock),
    .reset(sizeCounter_reset),
    .io_value_ready(sizeCounter_io_value_ready),
    .io_value_bits(sizeCounter_io_value_bits),
    .io_resetValue(sizeCounter_io_resetValue)
  );
  assign io_in_ready = sizeCounter_io_value_bits == io_in_bits_size & io_out_ready; // @[SizeHandler.scala 34:52 35:14 38:14]
  assign io_out_valid = io_in_valid; // @[SizeHandler.scala 25:16]
  assign io_out_bits_sel = io_in_bits_sel; // @[SizeHandler.scala 28:34]
  assign sizeCounter_clock = clock;
  assign sizeCounter_reset = reset;
  assign sizeCounter_io_value_ready = sizeCounter_io_value_bits == io_in_bits_size ? 1'h0 : fire; // @[SizeHandler.scala 34:52 Counter.scala 36:22 SizeHandler.scala 39:32]
  assign sizeCounter_io_resetValue = sizeCounter_io_value_bits == io_in_bits_size & fire; // @[SizeHandler.scala 34:52 Counter.scala 35:21 SizeHandler.scala 36:31]
endmodule
module Queue_26(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_sel,
  input  [13:0] io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_sel,
  output [13:0] io_deq_bits_size
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  ram_sel [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_sel_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_sel_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_sel_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_sel_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_sel_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_sel_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_sel_MPORT_en; // @[Decoupled.scala 259:95]
  reg [13:0] ram_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_10 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_10 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_sel_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sel_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_sel_io_deq_bits_MPORT_data = ram_sel[ram_sel_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_sel_MPORT_data = io_enq_bits_sel;
  assign ram_sel_MPORT_addr = 1'h0;
  assign ram_sel_MPORT_mask = 1'h1;
  assign ram_sel_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_sel = empty ? io_enq_bits_sel : ram_sel_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_sel_MPORT_en & ram_sel_MPORT_mask) begin
      ram_sel[ram_sel_MPORT_addr] <= ram_sel_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_sel[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[13:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_27(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_sel,
  input  [13:0] io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_sel,
  output [13:0] io_deq_bits_size
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  ram_sel [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_sel_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_sel_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_sel_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_sel_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_sel_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_sel_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_sel_MPORT_en; // @[Decoupled.scala 259:95]
  reg [13:0] ram_size [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [13:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [5:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [5:0] _value_T_1 = enq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire  _GEN_13 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_13 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire [5:0] _value_T_3 = deq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_sel_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sel_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_sel_io_deq_bits_MPORT_data = ram_sel[ram_sel_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_sel_MPORT_data = io_enq_bits_sel;
  assign ram_sel_MPORT_addr = enq_ptr_value;
  assign ram_sel_MPORT_mask = 1'h1;
  assign ram_sel_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_13 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | ~full; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_sel = empty ? io_enq_bits_sel : ram_sel_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_sel_MPORT_en & ram_sel_MPORT_mask) begin
      ram_sel[ram_sel_MPORT_addr] <= ram_sel_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_sel[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[13:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LocalRouter(
  input         clock,
  input         reset,
  output        io_control_ready,
  input         io_control_valid,
  input  [3:0]  io_control_bits_kind,
  input  [13:0] io_control_bits_size,
  output        io_mem_output_ready,
  input         io_mem_output_valid,
  input  [15:0] io_mem_output_bits_0,
  input  [15:0] io_mem_output_bits_1,
  input  [15:0] io_mem_output_bits_2,
  input  [15:0] io_mem_output_bits_3,
  input  [15:0] io_mem_output_bits_4,
  input  [15:0] io_mem_output_bits_5,
  input  [15:0] io_mem_output_bits_6,
  input  [15:0] io_mem_output_bits_7,
  input  [15:0] io_mem_output_bits_8,
  input  [15:0] io_mem_output_bits_9,
  input  [15:0] io_mem_output_bits_10,
  input  [15:0] io_mem_output_bits_11,
  input  [15:0] io_mem_output_bits_12,
  input  [15:0] io_mem_output_bits_13,
  input  [15:0] io_mem_output_bits_14,
  input  [15:0] io_mem_output_bits_15,
  input  [15:0] io_mem_output_bits_16,
  input  [15:0] io_mem_output_bits_17,
  input  [15:0] io_mem_output_bits_18,
  input  [15:0] io_mem_output_bits_19,
  input  [15:0] io_mem_output_bits_20,
  input  [15:0] io_mem_output_bits_21,
  input  [15:0] io_mem_output_bits_22,
  input  [15:0] io_mem_output_bits_23,
  input  [15:0] io_mem_output_bits_24,
  input  [15:0] io_mem_output_bits_25,
  input  [15:0] io_mem_output_bits_26,
  input  [15:0] io_mem_output_bits_27,
  input  [15:0] io_mem_output_bits_28,
  input  [15:0] io_mem_output_bits_29,
  input  [15:0] io_mem_output_bits_30,
  input  [15:0] io_mem_output_bits_31,
  input         io_mem_input_ready,
  output        io_mem_input_valid,
  output [15:0] io_mem_input_bits_0,
  output [15:0] io_mem_input_bits_1,
  output [15:0] io_mem_input_bits_2,
  output [15:0] io_mem_input_bits_3,
  output [15:0] io_mem_input_bits_4,
  output [15:0] io_mem_input_bits_5,
  output [15:0] io_mem_input_bits_6,
  output [15:0] io_mem_input_bits_7,
  output [15:0] io_mem_input_bits_8,
  output [15:0] io_mem_input_bits_9,
  output [15:0] io_mem_input_bits_10,
  output [15:0] io_mem_input_bits_11,
  output [15:0] io_mem_input_bits_12,
  output [15:0] io_mem_input_bits_13,
  output [15:0] io_mem_input_bits_14,
  output [15:0] io_mem_input_bits_15,
  output [15:0] io_mem_input_bits_16,
  output [15:0] io_mem_input_bits_17,
  output [15:0] io_mem_input_bits_18,
  output [15:0] io_mem_input_bits_19,
  output [15:0] io_mem_input_bits_20,
  output [15:0] io_mem_input_bits_21,
  output [15:0] io_mem_input_bits_22,
  output [15:0] io_mem_input_bits_23,
  output [15:0] io_mem_input_bits_24,
  output [15:0] io_mem_input_bits_25,
  output [15:0] io_mem_input_bits_26,
  output [15:0] io_mem_input_bits_27,
  output [15:0] io_mem_input_bits_28,
  output [15:0] io_mem_input_bits_29,
  output [15:0] io_mem_input_bits_30,
  output [15:0] io_mem_input_bits_31,
  input         io_array_input_ready,
  output        io_array_input_valid,
  output [15:0] io_array_input_bits_0,
  output [15:0] io_array_input_bits_1,
  output [15:0] io_array_input_bits_2,
  output [15:0] io_array_input_bits_3,
  output [15:0] io_array_input_bits_4,
  output [15:0] io_array_input_bits_5,
  output [15:0] io_array_input_bits_6,
  output [15:0] io_array_input_bits_7,
  output [15:0] io_array_input_bits_8,
  output [15:0] io_array_input_bits_9,
  output [15:0] io_array_input_bits_10,
  output [15:0] io_array_input_bits_11,
  output [15:0] io_array_input_bits_12,
  output [15:0] io_array_input_bits_13,
  output [15:0] io_array_input_bits_14,
  output [15:0] io_array_input_bits_15,
  output [15:0] io_array_input_bits_16,
  output [15:0] io_array_input_bits_17,
  output [15:0] io_array_input_bits_18,
  output [15:0] io_array_input_bits_19,
  output [15:0] io_array_input_bits_20,
  output [15:0] io_array_input_bits_21,
  output [15:0] io_array_input_bits_22,
  output [15:0] io_array_input_bits_23,
  output [15:0] io_array_input_bits_24,
  output [15:0] io_array_input_bits_25,
  output [15:0] io_array_input_bits_26,
  output [15:0] io_array_input_bits_27,
  output [15:0] io_array_input_bits_28,
  output [15:0] io_array_input_bits_29,
  output [15:0] io_array_input_bits_30,
  output [15:0] io_array_input_bits_31,
  output        io_array_output_ready,
  input         io_array_output_valid,
  input  [15:0] io_array_output_bits_0,
  input  [15:0] io_array_output_bits_1,
  input  [15:0] io_array_output_bits_2,
  input  [15:0] io_array_output_bits_3,
  input  [15:0] io_array_output_bits_4,
  input  [15:0] io_array_output_bits_5,
  input  [15:0] io_array_output_bits_6,
  input  [15:0] io_array_output_bits_7,
  input  [15:0] io_array_output_bits_8,
  input  [15:0] io_array_output_bits_9,
  input  [15:0] io_array_output_bits_10,
  input  [15:0] io_array_output_bits_11,
  input  [15:0] io_array_output_bits_12,
  input  [15:0] io_array_output_bits_13,
  input  [15:0] io_array_output_bits_14,
  input  [15:0] io_array_output_bits_15,
  input  [15:0] io_array_output_bits_16,
  input  [15:0] io_array_output_bits_17,
  input  [15:0] io_array_output_bits_18,
  input  [15:0] io_array_output_bits_19,
  input  [15:0] io_array_output_bits_20,
  input  [15:0] io_array_output_bits_21,
  input  [15:0] io_array_output_bits_22,
  input  [15:0] io_array_output_bits_23,
  input  [15:0] io_array_output_bits_24,
  input  [15:0] io_array_output_bits_25,
  input  [15:0] io_array_output_bits_26,
  input  [15:0] io_array_output_bits_27,
  input  [15:0] io_array_output_bits_28,
  input  [15:0] io_array_output_bits_29,
  input  [15:0] io_array_output_bits_30,
  input  [15:0] io_array_output_bits_31,
  input         io_array_weightInput_ready,
  output        io_array_weightInput_valid,
  output [15:0] io_array_weightInput_bits_0,
  output [15:0] io_array_weightInput_bits_1,
  output [15:0] io_array_weightInput_bits_2,
  output [15:0] io_array_weightInput_bits_3,
  output [15:0] io_array_weightInput_bits_4,
  output [15:0] io_array_weightInput_bits_5,
  output [15:0] io_array_weightInput_bits_6,
  output [15:0] io_array_weightInput_bits_7,
  output [15:0] io_array_weightInput_bits_8,
  output [15:0] io_array_weightInput_bits_9,
  output [15:0] io_array_weightInput_bits_10,
  output [15:0] io_array_weightInput_bits_11,
  output [15:0] io_array_weightInput_bits_12,
  output [15:0] io_array_weightInput_bits_13,
  output [15:0] io_array_weightInput_bits_14,
  output [15:0] io_array_weightInput_bits_15,
  output [15:0] io_array_weightInput_bits_16,
  output [15:0] io_array_weightInput_bits_17,
  output [15:0] io_array_weightInput_bits_18,
  output [15:0] io_array_weightInput_bits_19,
  output [15:0] io_array_weightInput_bits_20,
  output [15:0] io_array_weightInput_bits_21,
  output [15:0] io_array_weightInput_bits_22,
  output [15:0] io_array_weightInput_bits_23,
  output [15:0] io_array_weightInput_bits_24,
  output [15:0] io_array_weightInput_bits_25,
  output [15:0] io_array_weightInput_bits_26,
  output [15:0] io_array_weightInput_bits_27,
  output [15:0] io_array_weightInput_bits_28,
  output [15:0] io_array_weightInput_bits_29,
  output [15:0] io_array_weightInput_bits_30,
  output [15:0] io_array_weightInput_bits_31,
  output        io_acc_output_ready,
  input         io_acc_output_valid,
  input  [15:0] io_acc_output_bits_0,
  input  [15:0] io_acc_output_bits_1,
  input  [15:0] io_acc_output_bits_2,
  input  [15:0] io_acc_output_bits_3,
  input  [15:0] io_acc_output_bits_4,
  input  [15:0] io_acc_output_bits_5,
  input  [15:0] io_acc_output_bits_6,
  input  [15:0] io_acc_output_bits_7,
  input  [15:0] io_acc_output_bits_8,
  input  [15:0] io_acc_output_bits_9,
  input  [15:0] io_acc_output_bits_10,
  input  [15:0] io_acc_output_bits_11,
  input  [15:0] io_acc_output_bits_12,
  input  [15:0] io_acc_output_bits_13,
  input  [15:0] io_acc_output_bits_14,
  input  [15:0] io_acc_output_bits_15,
  input  [15:0] io_acc_output_bits_16,
  input  [15:0] io_acc_output_bits_17,
  input  [15:0] io_acc_output_bits_18,
  input  [15:0] io_acc_output_bits_19,
  input  [15:0] io_acc_output_bits_20,
  input  [15:0] io_acc_output_bits_21,
  input  [15:0] io_acc_output_bits_22,
  input  [15:0] io_acc_output_bits_23,
  input  [15:0] io_acc_output_bits_24,
  input  [15:0] io_acc_output_bits_25,
  input  [15:0] io_acc_output_bits_26,
  input  [15:0] io_acc_output_bits_27,
  input  [15:0] io_acc_output_bits_28,
  input  [15:0] io_acc_output_bits_29,
  input  [15:0] io_acc_output_bits_30,
  input  [15:0] io_acc_output_bits_31,
  input         io_acc_input_ready,
  output        io_acc_input_valid,
  output [15:0] io_acc_input_bits_0,
  output [15:0] io_acc_input_bits_1,
  output [15:0] io_acc_input_bits_2,
  output [15:0] io_acc_input_bits_3,
  output [15:0] io_acc_input_bits_4,
  output [15:0] io_acc_input_bits_5,
  output [15:0] io_acc_input_bits_6,
  output [15:0] io_acc_input_bits_7,
  output [15:0] io_acc_input_bits_8,
  output [15:0] io_acc_input_bits_9,
  output [15:0] io_acc_input_bits_10,
  output [15:0] io_acc_input_bits_11,
  output [15:0] io_acc_input_bits_12,
  output [15:0] io_acc_input_bits_13,
  output [15:0] io_acc_input_bits_14,
  output [15:0] io_acc_input_bits_15,
  output [15:0] io_acc_input_bits_16,
  output [15:0] io_acc_input_bits_17,
  output [15:0] io_acc_input_bits_18,
  output [15:0] io_acc_input_bits_19,
  output [15:0] io_acc_input_bits_20,
  output [15:0] io_acc_input_bits_21,
  output [15:0] io_acc_input_bits_22,
  output [15:0] io_acc_input_bits_23,
  output [15:0] io_acc_input_bits_24,
  output [15:0] io_acc_input_bits_25,
  output [15:0] io_acc_input_bits_26,
  output [15:0] io_acc_input_bits_27,
  output [15:0] io_acc_input_bits_28,
  output [15:0] io_acc_input_bits_29,
  output [15:0] io_acc_input_bits_30,
  output [15:0] io_acc_input_bits_31,
  input         io_timeout,
  input         io_tracepoint,
  input  [31:0] io_programCounter
);
  wire  memReadDataDemuxModule_io_in_ready; // @[LocalRouter.scala 55:38]
  wire  memReadDataDemuxModule_io_in_valid; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_0; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_1; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_2; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_3; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_4; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_5; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_6; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_7; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_8; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_9; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_10; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_11; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_12; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_13; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_14; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_15; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_16; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_17; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_18; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_19; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_20; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_21; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_22; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_23; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_24; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_25; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_26; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_27; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_28; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_29; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_30; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_in_bits_31; // @[LocalRouter.scala 55:38]
  wire  memReadDataDemuxModule_io_sel_ready; // @[LocalRouter.scala 55:38]
  wire  memReadDataDemuxModule_io_sel_valid; // @[LocalRouter.scala 55:38]
  wire [1:0] memReadDataDemuxModule_io_sel_bits; // @[LocalRouter.scala 55:38]
  wire  memReadDataDemuxModule_io_out_0_ready; // @[LocalRouter.scala 55:38]
  wire  memReadDataDemuxModule_io_out_0_valid; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_0; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_1; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_2; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_3; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_4; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_5; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_6; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_7; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_8; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_9; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_10; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_11; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_12; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_13; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_14; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_15; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_16; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_17; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_18; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_19; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_20; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_21; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_22; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_23; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_24; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_25; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_26; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_27; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_28; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_29; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_30; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_0_bits_31; // @[LocalRouter.scala 55:38]
  wire  memReadDataDemuxModule_io_out_1_ready; // @[LocalRouter.scala 55:38]
  wire  memReadDataDemuxModule_io_out_1_valid; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_0; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_1; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_2; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_3; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_4; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_5; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_6; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_7; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_8; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_9; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_10; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_11; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_12; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_13; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_14; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_15; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_16; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_17; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_18; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_19; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_20; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_21; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_22; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_23; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_24; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_25; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_26; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_27; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_28; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_29; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_30; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_1_bits_31; // @[LocalRouter.scala 55:38]
  wire  memReadDataDemuxModule_io_out_2_ready; // @[LocalRouter.scala 55:38]
  wire  memReadDataDemuxModule_io_out_2_valid; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_0; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_1; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_2; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_3; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_4; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_5; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_6; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_7; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_8; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_9; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_10; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_11; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_12; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_13; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_14; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_15; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_16; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_17; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_18; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_19; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_20; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_21; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_22; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_23; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_24; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_25; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_26; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_27; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_28; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_29; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_30; // @[LocalRouter.scala 55:38]
  wire [15:0] memReadDataDemuxModule_io_out_2_bits_31; // @[LocalRouter.scala 55:38]
  wire  memWriteDataMuxModule_io_in_0_ready; // @[LocalRouter.scala 66:37]
  wire  memWriteDataMuxModule_io_in_0_valid; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_0; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_1; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_2; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_3; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_4; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_5; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_6; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_7; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_8; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_9; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_10; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_11; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_12; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_13; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_14; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_15; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_16; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_17; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_18; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_19; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_20; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_21; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_22; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_23; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_24; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_25; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_26; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_27; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_28; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_29; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_30; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_0_bits_31; // @[LocalRouter.scala 66:37]
  wire  memWriteDataMuxModule_io_in_1_ready; // @[LocalRouter.scala 66:37]
  wire  memWriteDataMuxModule_io_in_1_valid; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_0; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_1; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_2; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_3; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_4; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_5; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_6; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_7; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_8; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_9; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_10; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_11; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_12; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_13; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_14; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_15; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_16; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_17; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_18; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_19; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_20; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_21; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_22; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_23; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_24; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_25; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_26; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_27; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_28; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_29; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_30; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_in_1_bits_31; // @[LocalRouter.scala 66:37]
  wire  memWriteDataMuxModule_io_sel_ready; // @[LocalRouter.scala 66:37]
  wire  memWriteDataMuxModule_io_sel_valid; // @[LocalRouter.scala 66:37]
  wire  memWriteDataMuxModule_io_sel_bits; // @[LocalRouter.scala 66:37]
  wire  memWriteDataMuxModule_io_out_ready; // @[LocalRouter.scala 66:37]
  wire  memWriteDataMuxModule_io_out_valid; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_0; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_1; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_2; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_3; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_4; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_5; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_6; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_7; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_8; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_9; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_10; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_11; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_12; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_13; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_14; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_15; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_16; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_17; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_18; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_19; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_20; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_21; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_22; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_23; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_24; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_25; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_26; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_27; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_28; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_29; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_30; // @[LocalRouter.scala 66:37]
  wire [15:0] memWriteDataMuxModule_io_out_bits_31; // @[LocalRouter.scala 66:37]
  wire  accWriteDataMuxModule_io_in_0_ready; // @[LocalRouter.scala 77:37]
  wire  accWriteDataMuxModule_io_in_0_valid; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_0; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_1; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_2; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_3; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_4; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_5; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_6; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_7; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_8; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_9; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_10; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_11; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_12; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_13; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_14; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_15; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_16; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_17; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_18; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_19; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_20; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_21; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_22; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_23; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_24; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_25; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_26; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_27; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_28; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_29; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_30; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_0_bits_31; // @[LocalRouter.scala 77:37]
  wire  accWriteDataMuxModule_io_in_1_ready; // @[LocalRouter.scala 77:37]
  wire  accWriteDataMuxModule_io_in_1_valid; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_0; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_1; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_2; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_3; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_4; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_5; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_6; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_7; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_8; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_9; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_10; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_11; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_12; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_13; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_14; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_15; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_16; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_17; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_18; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_19; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_20; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_21; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_22; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_23; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_24; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_25; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_26; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_27; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_28; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_29; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_30; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_in_1_bits_31; // @[LocalRouter.scala 77:37]
  wire  accWriteDataMuxModule_io_sel_ready; // @[LocalRouter.scala 77:37]
  wire  accWriteDataMuxModule_io_sel_valid; // @[LocalRouter.scala 77:37]
  wire  accWriteDataMuxModule_io_sel_bits; // @[LocalRouter.scala 77:37]
  wire  accWriteDataMuxModule_io_out_ready; // @[LocalRouter.scala 77:37]
  wire  accWriteDataMuxModule_io_out_valid; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_0; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_1; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_2; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_3; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_4; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_5; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_6; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_7; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_8; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_9; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_10; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_11; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_12; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_13; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_14; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_15; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_16; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_17; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_18; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_19; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_20; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_21; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_22; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_23; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_24; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_25; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_26; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_27; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_28; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_29; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_30; // @[LocalRouter.scala 77:37]
  wire [15:0] accWriteDataMuxModule_io_out_bits_31; // @[LocalRouter.scala 77:37]
  wire  sizeHandler_clock; // @[package.scala 33:29]
  wire  sizeHandler_reset; // @[package.scala 33:29]
  wire  sizeHandler_io_in_ready; // @[package.scala 33:29]
  wire  sizeHandler_io_in_valid; // @[package.scala 33:29]
  wire [1:0] sizeHandler_io_in_bits_sel; // @[package.scala 33:29]
  wire [13:0] sizeHandler_io_in_bits_size; // @[package.scala 33:29]
  wire  sizeHandler_io_out_ready; // @[package.scala 33:29]
  wire  sizeHandler_io_out_valid; // @[package.scala 33:29]
  wire [1:0] sizeHandler_io_out_bits_sel; // @[package.scala 33:29]
  wire  memReadDataDemux_clock; // @[Mem.scala 22:19]
  wire  memReadDataDemux_reset; // @[Mem.scala 22:19]
  wire  memReadDataDemux_io_enq_ready; // @[Mem.scala 22:19]
  wire  memReadDataDemux_io_enq_valid; // @[Mem.scala 22:19]
  wire [1:0] memReadDataDemux_io_enq_bits_sel; // @[Mem.scala 22:19]
  wire [13:0] memReadDataDemux_io_enq_bits_size; // @[Mem.scala 22:19]
  wire  memReadDataDemux_io_deq_ready; // @[Mem.scala 22:19]
  wire  memReadDataDemux_io_deq_valid; // @[Mem.scala 22:19]
  wire [1:0] memReadDataDemux_io_deq_bits_sel; // @[Mem.scala 22:19]
  wire [13:0] memReadDataDemux_io_deq_bits_size; // @[Mem.scala 22:19]
  wire  sizeHandler_1_clock; // @[package.scala 33:29]
  wire  sizeHandler_1_reset; // @[package.scala 33:29]
  wire  sizeHandler_1_io_in_ready; // @[package.scala 33:29]
  wire  sizeHandler_1_io_in_valid; // @[package.scala 33:29]
  wire  sizeHandler_1_io_in_bits_sel; // @[package.scala 33:29]
  wire [13:0] sizeHandler_1_io_in_bits_size; // @[package.scala 33:29]
  wire  sizeHandler_1_io_out_ready; // @[package.scala 33:29]
  wire  sizeHandler_1_io_out_valid; // @[package.scala 33:29]
  wire  sizeHandler_1_io_out_bits_sel; // @[package.scala 33:29]
  wire  memWriteDataMux_clock; // @[Mem.scala 22:19]
  wire  memWriteDataMux_reset; // @[Mem.scala 22:19]
  wire  memWriteDataMux_io_enq_ready; // @[Mem.scala 22:19]
  wire  memWriteDataMux_io_enq_valid; // @[Mem.scala 22:19]
  wire  memWriteDataMux_io_enq_bits_sel; // @[Mem.scala 22:19]
  wire [13:0] memWriteDataMux_io_enq_bits_size; // @[Mem.scala 22:19]
  wire  memWriteDataMux_io_deq_ready; // @[Mem.scala 22:19]
  wire  memWriteDataMux_io_deq_valid; // @[Mem.scala 22:19]
  wire  memWriteDataMux_io_deq_bits_sel; // @[Mem.scala 22:19]
  wire [13:0] memWriteDataMux_io_deq_bits_size; // @[Mem.scala 22:19]
  wire  sizeHandler_2_clock; // @[package.scala 33:29]
  wire  sizeHandler_2_reset; // @[package.scala 33:29]
  wire  sizeHandler_2_io_in_ready; // @[package.scala 33:29]
  wire  sizeHandler_2_io_in_valid; // @[package.scala 33:29]
  wire  sizeHandler_2_io_in_bits_sel; // @[package.scala 33:29]
  wire [13:0] sizeHandler_2_io_in_bits_size; // @[package.scala 33:29]
  wire  sizeHandler_2_io_out_ready; // @[package.scala 33:29]
  wire  sizeHandler_2_io_out_valid; // @[package.scala 33:29]
  wire  sizeHandler_2_io_out_bits_sel; // @[package.scala 33:29]
  wire  accWriteDataMux_clock; // @[Mem.scala 22:19]
  wire  accWriteDataMux_reset; // @[Mem.scala 22:19]
  wire  accWriteDataMux_io_enq_ready; // @[Mem.scala 22:19]
  wire  accWriteDataMux_io_enq_valid; // @[Mem.scala 22:19]
  wire  accWriteDataMux_io_enq_bits_sel; // @[Mem.scala 22:19]
  wire [13:0] accWriteDataMux_io_enq_bits_size; // @[Mem.scala 22:19]
  wire  accWriteDataMux_io_deq_ready; // @[Mem.scala 22:19]
  wire  accWriteDataMux_io_deq_valid; // @[Mem.scala 22:19]
  wire  accWriteDataMux_io_deq_bits_sel; // @[Mem.scala 22:19]
  wire [13:0] accWriteDataMux_io_deq_bits_size; // @[Mem.scala 22:19]
  wire  enqueuer1_clock; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer1_reset; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer1_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer1_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer1_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer1_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_clock; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_reset; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  enqueuer2_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  _T_3 = io_control_bits_kind == 4'h4; // @[LocalRouter.scala 143:32]
  wire  _T_4 = io_control_bits_kind == 4'h5; // @[LocalRouter.scala 150:23]
  wire  _GEN_0 = _T_4 & io_control_valid; // @[LocalRouter.scala 151:5 MultiEnqueue.scala 40:17 84:17]
  wire  io_control_ready_memReadDataDemux_io_enq_w_2_ready = memReadDataDemux_io_enq_ready; // @[ReadyValid.scala 16:17 MultiEnqueue.scala 85:10]
  wire  _GEN_1 = _T_4 & io_control_ready_memReadDataDemux_io_enq_w_2_ready; // @[LocalRouter.scala 151:5 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  io_control_ready_memReadDataDemux_io_enq_w_2_valid = enqueuer2_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_2 = _T_4 & io_control_ready_memReadDataDemux_io_enq_w_2_valid; // @[LocalRouter.scala 151:5 MultiEnqueue.scala 85:10 package.scala 405:15]
  wire [1:0] _GEN_3 = _T_4 ? 2'h2 : 2'h0; // @[LocalRouter.scala 151:5 MultiEnqueue.scala 85:10 package.scala 404:14]
  wire [13:0] _GEN_4 = _T_4 ? io_control_bits_size : 14'h0; // @[LocalRouter.scala 151:5 MultiEnqueue.scala 85:10 package.scala 404:14]
  wire  io_control_ready_accWriteDataMux_io_enq_w_2_ready = accWriteDataMux_io_enq_ready; // @[ReadyValid.scala 16:17 MultiEnqueue.scala 86:10]
  wire  _GEN_5 = _T_4 & io_control_ready_accWriteDataMux_io_enq_w_2_ready; // @[LocalRouter.scala 151:5 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  io_control_ready_accWriteDataMux_io_enq_w_2_valid = enqueuer2_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_6 = _T_4 & io_control_ready_accWriteDataMux_io_enq_w_2_valid; // @[LocalRouter.scala 151:5 MultiEnqueue.scala 86:10 package.scala 405:15]
  wire  _GEN_9 = _T_4 ? enqueuer2_io_in_ready : 1'h1; // @[LocalRouter.scala 151:5 152:19 160:19]
  wire  _GEN_10 = io_control_bits_kind == 4'h4 & io_control_valid; // @[LocalRouter.scala 143:78 MultiEnqueue.scala 40:17 60:17]
  wire  io_control_ready_memWriteDataMux_io_enq_w_ready = memWriteDataMux_io_enq_ready; // @[ReadyValid.scala 16:17 MultiEnqueue.scala 61:10]
  wire  _GEN_11 = io_control_bits_kind == 4'h4 & io_control_ready_memWriteDataMux_io_enq_w_ready; // @[LocalRouter.scala 143:78 ReadyValid.scala 19:11 MultiEnqueue.scala 42:18]
  wire  io_control_ready_memWriteDataMux_io_enq_w_valid = enqueuer1_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_12 = io_control_bits_kind == 4'h4 & io_control_ready_memWriteDataMux_io_enq_w_valid; // @[LocalRouter.scala 143:78 MultiEnqueue.scala 61:10 package.scala 405:15]
  wire [13:0] _GEN_14 = io_control_bits_kind == 4'h4 ? io_control_bits_size : 14'h0; // @[LocalRouter.scala 143:78 MultiEnqueue.scala 61:10 package.scala 404:14]
  wire  _GEN_15 = io_control_bits_kind == 4'h4 ? enqueuer1_io_in_ready : _GEN_9; // @[LocalRouter.scala 143:78 144:19]
  wire  _GEN_16 = io_control_bits_kind == 4'h4 ? 1'h0 : _GEN_0; // @[LocalRouter.scala 143:78 MultiEnqueue.scala 40:17]
  wire  _GEN_17 = io_control_bits_kind == 4'h4 ? 1'h0 : _GEN_1; // @[LocalRouter.scala 143:78 MultiEnqueue.scala 42:18]
  wire  _GEN_18 = io_control_bits_kind == 4'h4 ? 1'h0 : _GEN_2; // @[LocalRouter.scala 143:78 package.scala 405:15]
  wire [1:0] _GEN_19 = io_control_bits_kind == 4'h4 ? 2'h0 : _GEN_3; // @[LocalRouter.scala 143:78 package.scala 404:14]
  wire [13:0] _GEN_20 = io_control_bits_kind == 4'h4 ? 14'h0 : _GEN_4; // @[LocalRouter.scala 143:78 package.scala 404:14]
  wire  _GEN_21 = io_control_bits_kind == 4'h4 ? 1'h0 : _GEN_5; // @[LocalRouter.scala 143:78 MultiEnqueue.scala 42:18]
  wire  _GEN_22 = io_control_bits_kind == 4'h4 ? 1'h0 : _GEN_6; // @[LocalRouter.scala 143:78 package.scala 405:15]
  wire  _GEN_23 = io_control_bits_kind == 4'h4 ? 1'h0 : _T_4; // @[LocalRouter.scala 143:78 package.scala 404:14]
  wire  _GEN_25 = io_control_bits_kind == 4'h3 ? io_control_valid : _GEN_10; // @[LocalRouter.scala 137:70 MultiEnqueue.scala 60:17]
  wire  _GEN_26 = io_control_bits_kind == 4'h3 ? io_control_ready_accWriteDataMux_io_enq_w_2_ready : _GEN_11; // @[LocalRouter.scala 137:70 ReadyValid.scala 19:11]
  wire  _GEN_27 = io_control_bits_kind == 4'h3 ? io_control_ready_memWriteDataMux_io_enq_w_valid : _GEN_22; // @[LocalRouter.scala 137:70 MultiEnqueue.scala 61:10]
  wire  _GEN_28 = io_control_bits_kind == 4'h3 ? 1'h0 : _GEN_23; // @[LocalRouter.scala 137:70 MultiEnqueue.scala 61:10]
  wire [13:0] _GEN_29 = io_control_bits_kind == 4'h3 ? io_control_bits_size : _GEN_20; // @[LocalRouter.scala 137:70 MultiEnqueue.scala 61:10]
  wire  _GEN_30 = io_control_bits_kind == 4'h3 ? enqueuer1_io_in_ready : _GEN_15; // @[LocalRouter.scala 137:70 138:19]
  wire  _GEN_31 = io_control_bits_kind == 4'h3 ? 1'h0 : _GEN_12; // @[LocalRouter.scala 137:70 package.scala 405:15]
  wire  _GEN_32 = io_control_bits_kind == 4'h3 ? 1'h0 : _T_3; // @[LocalRouter.scala 137:70 package.scala 404:14]
  wire [13:0] _GEN_33 = io_control_bits_kind == 4'h3 ? 14'h0 : _GEN_14; // @[LocalRouter.scala 137:70 package.scala 404:14]
  wire  _GEN_34 = io_control_bits_kind == 4'h3 ? 1'h0 : _GEN_16; // @[LocalRouter.scala 137:70 MultiEnqueue.scala 40:17]
  wire  _GEN_35 = io_control_bits_kind == 4'h3 ? 1'h0 : _GEN_17; // @[LocalRouter.scala 137:70 MultiEnqueue.scala 42:18]
  wire  _GEN_36 = io_control_bits_kind == 4'h3 ? 1'h0 : _GEN_18; // @[LocalRouter.scala 137:70 package.scala 405:15]
  wire [1:0] _GEN_37 = io_control_bits_kind == 4'h3 ? 2'h0 : _GEN_19; // @[LocalRouter.scala 137:70 package.scala 404:14]
  wire [13:0] _GEN_38 = io_control_bits_kind == 4'h3 ? 14'h0 : _GEN_20; // @[LocalRouter.scala 137:70 package.scala 404:14]
  wire  _GEN_39 = io_control_bits_kind == 4'h3 ? 1'h0 : _GEN_21; // @[LocalRouter.scala 137:70 MultiEnqueue.scala 42:18]
  wire  _GEN_40 = io_control_bits_kind == 4'h2 ? io_control_valid : _GEN_34; // @[LocalRouter.scala 129:78 MultiEnqueue.scala 84:17]
  wire  _GEN_41 = io_control_bits_kind == 4'h2 ? io_control_ready_memReadDataDemux_io_enq_w_2_ready : _GEN_35; // @[LocalRouter.scala 129:78 ReadyValid.scala 19:11]
  wire  _GEN_42 = io_control_bits_kind == 4'h2 ? io_control_ready_memReadDataDemux_io_enq_w_2_valid : _GEN_36; // @[LocalRouter.scala 129:78 MultiEnqueue.scala 85:10]
  wire [1:0] _GEN_43 = io_control_bits_kind == 4'h2 ? 2'h1 : _GEN_37; // @[LocalRouter.scala 129:78 MultiEnqueue.scala 85:10]
  wire [13:0] _GEN_44 = io_control_bits_kind == 4'h2 ? io_control_bits_size : _GEN_38; // @[LocalRouter.scala 129:78 MultiEnqueue.scala 85:10]
  wire  _GEN_45 = io_control_bits_kind == 4'h2 ? io_control_ready_accWriteDataMux_io_enq_w_2_ready : _GEN_39; // @[LocalRouter.scala 129:78 ReadyValid.scala 19:11]
  wire  _GEN_46 = io_control_bits_kind == 4'h2 ? io_control_ready_accWriteDataMux_io_enq_w_2_valid : _GEN_27; // @[LocalRouter.scala 129:78 MultiEnqueue.scala 86:10]
  wire  _GEN_47 = io_control_bits_kind == 4'h2 ? 1'h0 : _GEN_28; // @[LocalRouter.scala 129:78 MultiEnqueue.scala 86:10]
  wire [13:0] _GEN_48 = io_control_bits_kind == 4'h2 ? io_control_bits_size : _GEN_29; // @[LocalRouter.scala 129:78 MultiEnqueue.scala 86:10]
  wire  _GEN_49 = io_control_bits_kind == 4'h2 ? enqueuer2_io_in_ready : _GEN_30; // @[LocalRouter.scala 129:78 130:19]
  wire  _GEN_50 = io_control_bits_kind == 4'h2 ? 1'h0 : _GEN_25; // @[LocalRouter.scala 129:78 MultiEnqueue.scala 40:17]
  wire  _GEN_51 = io_control_bits_kind == 4'h2 ? 1'h0 : _GEN_26; // @[LocalRouter.scala 129:78 MultiEnqueue.scala 42:18]
  wire  _GEN_52 = io_control_bits_kind == 4'h2 ? 1'h0 : _GEN_31; // @[LocalRouter.scala 129:78 package.scala 405:15]
  wire  _GEN_53 = io_control_bits_kind == 4'h2 ? 1'h0 : _GEN_32; // @[LocalRouter.scala 129:78 package.scala 404:14]
  wire [13:0] _GEN_54 = io_control_bits_kind == 4'h2 ? 14'h0 : _GEN_33; // @[LocalRouter.scala 129:78 package.scala 404:14]
  Demux_3 memReadDataDemuxModule ( // @[LocalRouter.scala 55:38]
    .io_in_ready(memReadDataDemuxModule_io_in_ready),
    .io_in_valid(memReadDataDemuxModule_io_in_valid),
    .io_in_bits_0(memReadDataDemuxModule_io_in_bits_0),
    .io_in_bits_1(memReadDataDemuxModule_io_in_bits_1),
    .io_in_bits_2(memReadDataDemuxModule_io_in_bits_2),
    .io_in_bits_3(memReadDataDemuxModule_io_in_bits_3),
    .io_in_bits_4(memReadDataDemuxModule_io_in_bits_4),
    .io_in_bits_5(memReadDataDemuxModule_io_in_bits_5),
    .io_in_bits_6(memReadDataDemuxModule_io_in_bits_6),
    .io_in_bits_7(memReadDataDemuxModule_io_in_bits_7),
    .io_in_bits_8(memReadDataDemuxModule_io_in_bits_8),
    .io_in_bits_9(memReadDataDemuxModule_io_in_bits_9),
    .io_in_bits_10(memReadDataDemuxModule_io_in_bits_10),
    .io_in_bits_11(memReadDataDemuxModule_io_in_bits_11),
    .io_in_bits_12(memReadDataDemuxModule_io_in_bits_12),
    .io_in_bits_13(memReadDataDemuxModule_io_in_bits_13),
    .io_in_bits_14(memReadDataDemuxModule_io_in_bits_14),
    .io_in_bits_15(memReadDataDemuxModule_io_in_bits_15),
    .io_in_bits_16(memReadDataDemuxModule_io_in_bits_16),
    .io_in_bits_17(memReadDataDemuxModule_io_in_bits_17),
    .io_in_bits_18(memReadDataDemuxModule_io_in_bits_18),
    .io_in_bits_19(memReadDataDemuxModule_io_in_bits_19),
    .io_in_bits_20(memReadDataDemuxModule_io_in_bits_20),
    .io_in_bits_21(memReadDataDemuxModule_io_in_bits_21),
    .io_in_bits_22(memReadDataDemuxModule_io_in_bits_22),
    .io_in_bits_23(memReadDataDemuxModule_io_in_bits_23),
    .io_in_bits_24(memReadDataDemuxModule_io_in_bits_24),
    .io_in_bits_25(memReadDataDemuxModule_io_in_bits_25),
    .io_in_bits_26(memReadDataDemuxModule_io_in_bits_26),
    .io_in_bits_27(memReadDataDemuxModule_io_in_bits_27),
    .io_in_bits_28(memReadDataDemuxModule_io_in_bits_28),
    .io_in_bits_29(memReadDataDemuxModule_io_in_bits_29),
    .io_in_bits_30(memReadDataDemuxModule_io_in_bits_30),
    .io_in_bits_31(memReadDataDemuxModule_io_in_bits_31),
    .io_sel_ready(memReadDataDemuxModule_io_sel_ready),
    .io_sel_valid(memReadDataDemuxModule_io_sel_valid),
    .io_sel_bits(memReadDataDemuxModule_io_sel_bits),
    .io_out_0_ready(memReadDataDemuxModule_io_out_0_ready),
    .io_out_0_valid(memReadDataDemuxModule_io_out_0_valid),
    .io_out_0_bits_0(memReadDataDemuxModule_io_out_0_bits_0),
    .io_out_0_bits_1(memReadDataDemuxModule_io_out_0_bits_1),
    .io_out_0_bits_2(memReadDataDemuxModule_io_out_0_bits_2),
    .io_out_0_bits_3(memReadDataDemuxModule_io_out_0_bits_3),
    .io_out_0_bits_4(memReadDataDemuxModule_io_out_0_bits_4),
    .io_out_0_bits_5(memReadDataDemuxModule_io_out_0_bits_5),
    .io_out_0_bits_6(memReadDataDemuxModule_io_out_0_bits_6),
    .io_out_0_bits_7(memReadDataDemuxModule_io_out_0_bits_7),
    .io_out_0_bits_8(memReadDataDemuxModule_io_out_0_bits_8),
    .io_out_0_bits_9(memReadDataDemuxModule_io_out_0_bits_9),
    .io_out_0_bits_10(memReadDataDemuxModule_io_out_0_bits_10),
    .io_out_0_bits_11(memReadDataDemuxModule_io_out_0_bits_11),
    .io_out_0_bits_12(memReadDataDemuxModule_io_out_0_bits_12),
    .io_out_0_bits_13(memReadDataDemuxModule_io_out_0_bits_13),
    .io_out_0_bits_14(memReadDataDemuxModule_io_out_0_bits_14),
    .io_out_0_bits_15(memReadDataDemuxModule_io_out_0_bits_15),
    .io_out_0_bits_16(memReadDataDemuxModule_io_out_0_bits_16),
    .io_out_0_bits_17(memReadDataDemuxModule_io_out_0_bits_17),
    .io_out_0_bits_18(memReadDataDemuxModule_io_out_0_bits_18),
    .io_out_0_bits_19(memReadDataDemuxModule_io_out_0_bits_19),
    .io_out_0_bits_20(memReadDataDemuxModule_io_out_0_bits_20),
    .io_out_0_bits_21(memReadDataDemuxModule_io_out_0_bits_21),
    .io_out_0_bits_22(memReadDataDemuxModule_io_out_0_bits_22),
    .io_out_0_bits_23(memReadDataDemuxModule_io_out_0_bits_23),
    .io_out_0_bits_24(memReadDataDemuxModule_io_out_0_bits_24),
    .io_out_0_bits_25(memReadDataDemuxModule_io_out_0_bits_25),
    .io_out_0_bits_26(memReadDataDemuxModule_io_out_0_bits_26),
    .io_out_0_bits_27(memReadDataDemuxModule_io_out_0_bits_27),
    .io_out_0_bits_28(memReadDataDemuxModule_io_out_0_bits_28),
    .io_out_0_bits_29(memReadDataDemuxModule_io_out_0_bits_29),
    .io_out_0_bits_30(memReadDataDemuxModule_io_out_0_bits_30),
    .io_out_0_bits_31(memReadDataDemuxModule_io_out_0_bits_31),
    .io_out_1_ready(memReadDataDemuxModule_io_out_1_ready),
    .io_out_1_valid(memReadDataDemuxModule_io_out_1_valid),
    .io_out_1_bits_0(memReadDataDemuxModule_io_out_1_bits_0),
    .io_out_1_bits_1(memReadDataDemuxModule_io_out_1_bits_1),
    .io_out_1_bits_2(memReadDataDemuxModule_io_out_1_bits_2),
    .io_out_1_bits_3(memReadDataDemuxModule_io_out_1_bits_3),
    .io_out_1_bits_4(memReadDataDemuxModule_io_out_1_bits_4),
    .io_out_1_bits_5(memReadDataDemuxModule_io_out_1_bits_5),
    .io_out_1_bits_6(memReadDataDemuxModule_io_out_1_bits_6),
    .io_out_1_bits_7(memReadDataDemuxModule_io_out_1_bits_7),
    .io_out_1_bits_8(memReadDataDemuxModule_io_out_1_bits_8),
    .io_out_1_bits_9(memReadDataDemuxModule_io_out_1_bits_9),
    .io_out_1_bits_10(memReadDataDemuxModule_io_out_1_bits_10),
    .io_out_1_bits_11(memReadDataDemuxModule_io_out_1_bits_11),
    .io_out_1_bits_12(memReadDataDemuxModule_io_out_1_bits_12),
    .io_out_1_bits_13(memReadDataDemuxModule_io_out_1_bits_13),
    .io_out_1_bits_14(memReadDataDemuxModule_io_out_1_bits_14),
    .io_out_1_bits_15(memReadDataDemuxModule_io_out_1_bits_15),
    .io_out_1_bits_16(memReadDataDemuxModule_io_out_1_bits_16),
    .io_out_1_bits_17(memReadDataDemuxModule_io_out_1_bits_17),
    .io_out_1_bits_18(memReadDataDemuxModule_io_out_1_bits_18),
    .io_out_1_bits_19(memReadDataDemuxModule_io_out_1_bits_19),
    .io_out_1_bits_20(memReadDataDemuxModule_io_out_1_bits_20),
    .io_out_1_bits_21(memReadDataDemuxModule_io_out_1_bits_21),
    .io_out_1_bits_22(memReadDataDemuxModule_io_out_1_bits_22),
    .io_out_1_bits_23(memReadDataDemuxModule_io_out_1_bits_23),
    .io_out_1_bits_24(memReadDataDemuxModule_io_out_1_bits_24),
    .io_out_1_bits_25(memReadDataDemuxModule_io_out_1_bits_25),
    .io_out_1_bits_26(memReadDataDemuxModule_io_out_1_bits_26),
    .io_out_1_bits_27(memReadDataDemuxModule_io_out_1_bits_27),
    .io_out_1_bits_28(memReadDataDemuxModule_io_out_1_bits_28),
    .io_out_1_bits_29(memReadDataDemuxModule_io_out_1_bits_29),
    .io_out_1_bits_30(memReadDataDemuxModule_io_out_1_bits_30),
    .io_out_1_bits_31(memReadDataDemuxModule_io_out_1_bits_31),
    .io_out_2_ready(memReadDataDemuxModule_io_out_2_ready),
    .io_out_2_valid(memReadDataDemuxModule_io_out_2_valid),
    .io_out_2_bits_0(memReadDataDemuxModule_io_out_2_bits_0),
    .io_out_2_bits_1(memReadDataDemuxModule_io_out_2_bits_1),
    .io_out_2_bits_2(memReadDataDemuxModule_io_out_2_bits_2),
    .io_out_2_bits_3(memReadDataDemuxModule_io_out_2_bits_3),
    .io_out_2_bits_4(memReadDataDemuxModule_io_out_2_bits_4),
    .io_out_2_bits_5(memReadDataDemuxModule_io_out_2_bits_5),
    .io_out_2_bits_6(memReadDataDemuxModule_io_out_2_bits_6),
    .io_out_2_bits_7(memReadDataDemuxModule_io_out_2_bits_7),
    .io_out_2_bits_8(memReadDataDemuxModule_io_out_2_bits_8),
    .io_out_2_bits_9(memReadDataDemuxModule_io_out_2_bits_9),
    .io_out_2_bits_10(memReadDataDemuxModule_io_out_2_bits_10),
    .io_out_2_bits_11(memReadDataDemuxModule_io_out_2_bits_11),
    .io_out_2_bits_12(memReadDataDemuxModule_io_out_2_bits_12),
    .io_out_2_bits_13(memReadDataDemuxModule_io_out_2_bits_13),
    .io_out_2_bits_14(memReadDataDemuxModule_io_out_2_bits_14),
    .io_out_2_bits_15(memReadDataDemuxModule_io_out_2_bits_15),
    .io_out_2_bits_16(memReadDataDemuxModule_io_out_2_bits_16),
    .io_out_2_bits_17(memReadDataDemuxModule_io_out_2_bits_17),
    .io_out_2_bits_18(memReadDataDemuxModule_io_out_2_bits_18),
    .io_out_2_bits_19(memReadDataDemuxModule_io_out_2_bits_19),
    .io_out_2_bits_20(memReadDataDemuxModule_io_out_2_bits_20),
    .io_out_2_bits_21(memReadDataDemuxModule_io_out_2_bits_21),
    .io_out_2_bits_22(memReadDataDemuxModule_io_out_2_bits_22),
    .io_out_2_bits_23(memReadDataDemuxModule_io_out_2_bits_23),
    .io_out_2_bits_24(memReadDataDemuxModule_io_out_2_bits_24),
    .io_out_2_bits_25(memReadDataDemuxModule_io_out_2_bits_25),
    .io_out_2_bits_26(memReadDataDemuxModule_io_out_2_bits_26),
    .io_out_2_bits_27(memReadDataDemuxModule_io_out_2_bits_27),
    .io_out_2_bits_28(memReadDataDemuxModule_io_out_2_bits_28),
    .io_out_2_bits_29(memReadDataDemuxModule_io_out_2_bits_29),
    .io_out_2_bits_30(memReadDataDemuxModule_io_out_2_bits_30),
    .io_out_2_bits_31(memReadDataDemuxModule_io_out_2_bits_31)
  );
  Mux memWriteDataMuxModule ( // @[LocalRouter.scala 66:37]
    .io_in_0_ready(memWriteDataMuxModule_io_in_0_ready),
    .io_in_0_valid(memWriteDataMuxModule_io_in_0_valid),
    .io_in_0_bits_0(memWriteDataMuxModule_io_in_0_bits_0),
    .io_in_0_bits_1(memWriteDataMuxModule_io_in_0_bits_1),
    .io_in_0_bits_2(memWriteDataMuxModule_io_in_0_bits_2),
    .io_in_0_bits_3(memWriteDataMuxModule_io_in_0_bits_3),
    .io_in_0_bits_4(memWriteDataMuxModule_io_in_0_bits_4),
    .io_in_0_bits_5(memWriteDataMuxModule_io_in_0_bits_5),
    .io_in_0_bits_6(memWriteDataMuxModule_io_in_0_bits_6),
    .io_in_0_bits_7(memWriteDataMuxModule_io_in_0_bits_7),
    .io_in_0_bits_8(memWriteDataMuxModule_io_in_0_bits_8),
    .io_in_0_bits_9(memWriteDataMuxModule_io_in_0_bits_9),
    .io_in_0_bits_10(memWriteDataMuxModule_io_in_0_bits_10),
    .io_in_0_bits_11(memWriteDataMuxModule_io_in_0_bits_11),
    .io_in_0_bits_12(memWriteDataMuxModule_io_in_0_bits_12),
    .io_in_0_bits_13(memWriteDataMuxModule_io_in_0_bits_13),
    .io_in_0_bits_14(memWriteDataMuxModule_io_in_0_bits_14),
    .io_in_0_bits_15(memWriteDataMuxModule_io_in_0_bits_15),
    .io_in_0_bits_16(memWriteDataMuxModule_io_in_0_bits_16),
    .io_in_0_bits_17(memWriteDataMuxModule_io_in_0_bits_17),
    .io_in_0_bits_18(memWriteDataMuxModule_io_in_0_bits_18),
    .io_in_0_bits_19(memWriteDataMuxModule_io_in_0_bits_19),
    .io_in_0_bits_20(memWriteDataMuxModule_io_in_0_bits_20),
    .io_in_0_bits_21(memWriteDataMuxModule_io_in_0_bits_21),
    .io_in_0_bits_22(memWriteDataMuxModule_io_in_0_bits_22),
    .io_in_0_bits_23(memWriteDataMuxModule_io_in_0_bits_23),
    .io_in_0_bits_24(memWriteDataMuxModule_io_in_0_bits_24),
    .io_in_0_bits_25(memWriteDataMuxModule_io_in_0_bits_25),
    .io_in_0_bits_26(memWriteDataMuxModule_io_in_0_bits_26),
    .io_in_0_bits_27(memWriteDataMuxModule_io_in_0_bits_27),
    .io_in_0_bits_28(memWriteDataMuxModule_io_in_0_bits_28),
    .io_in_0_bits_29(memWriteDataMuxModule_io_in_0_bits_29),
    .io_in_0_bits_30(memWriteDataMuxModule_io_in_0_bits_30),
    .io_in_0_bits_31(memWriteDataMuxModule_io_in_0_bits_31),
    .io_in_1_ready(memWriteDataMuxModule_io_in_1_ready),
    .io_in_1_valid(memWriteDataMuxModule_io_in_1_valid),
    .io_in_1_bits_0(memWriteDataMuxModule_io_in_1_bits_0),
    .io_in_1_bits_1(memWriteDataMuxModule_io_in_1_bits_1),
    .io_in_1_bits_2(memWriteDataMuxModule_io_in_1_bits_2),
    .io_in_1_bits_3(memWriteDataMuxModule_io_in_1_bits_3),
    .io_in_1_bits_4(memWriteDataMuxModule_io_in_1_bits_4),
    .io_in_1_bits_5(memWriteDataMuxModule_io_in_1_bits_5),
    .io_in_1_bits_6(memWriteDataMuxModule_io_in_1_bits_6),
    .io_in_1_bits_7(memWriteDataMuxModule_io_in_1_bits_7),
    .io_in_1_bits_8(memWriteDataMuxModule_io_in_1_bits_8),
    .io_in_1_bits_9(memWriteDataMuxModule_io_in_1_bits_9),
    .io_in_1_bits_10(memWriteDataMuxModule_io_in_1_bits_10),
    .io_in_1_bits_11(memWriteDataMuxModule_io_in_1_bits_11),
    .io_in_1_bits_12(memWriteDataMuxModule_io_in_1_bits_12),
    .io_in_1_bits_13(memWriteDataMuxModule_io_in_1_bits_13),
    .io_in_1_bits_14(memWriteDataMuxModule_io_in_1_bits_14),
    .io_in_1_bits_15(memWriteDataMuxModule_io_in_1_bits_15),
    .io_in_1_bits_16(memWriteDataMuxModule_io_in_1_bits_16),
    .io_in_1_bits_17(memWriteDataMuxModule_io_in_1_bits_17),
    .io_in_1_bits_18(memWriteDataMuxModule_io_in_1_bits_18),
    .io_in_1_bits_19(memWriteDataMuxModule_io_in_1_bits_19),
    .io_in_1_bits_20(memWriteDataMuxModule_io_in_1_bits_20),
    .io_in_1_bits_21(memWriteDataMuxModule_io_in_1_bits_21),
    .io_in_1_bits_22(memWriteDataMuxModule_io_in_1_bits_22),
    .io_in_1_bits_23(memWriteDataMuxModule_io_in_1_bits_23),
    .io_in_1_bits_24(memWriteDataMuxModule_io_in_1_bits_24),
    .io_in_1_bits_25(memWriteDataMuxModule_io_in_1_bits_25),
    .io_in_1_bits_26(memWriteDataMuxModule_io_in_1_bits_26),
    .io_in_1_bits_27(memWriteDataMuxModule_io_in_1_bits_27),
    .io_in_1_bits_28(memWriteDataMuxModule_io_in_1_bits_28),
    .io_in_1_bits_29(memWriteDataMuxModule_io_in_1_bits_29),
    .io_in_1_bits_30(memWriteDataMuxModule_io_in_1_bits_30),
    .io_in_1_bits_31(memWriteDataMuxModule_io_in_1_bits_31),
    .io_sel_ready(memWriteDataMuxModule_io_sel_ready),
    .io_sel_valid(memWriteDataMuxModule_io_sel_valid),
    .io_sel_bits(memWriteDataMuxModule_io_sel_bits),
    .io_out_ready(memWriteDataMuxModule_io_out_ready),
    .io_out_valid(memWriteDataMuxModule_io_out_valid),
    .io_out_bits_0(memWriteDataMuxModule_io_out_bits_0),
    .io_out_bits_1(memWriteDataMuxModule_io_out_bits_1),
    .io_out_bits_2(memWriteDataMuxModule_io_out_bits_2),
    .io_out_bits_3(memWriteDataMuxModule_io_out_bits_3),
    .io_out_bits_4(memWriteDataMuxModule_io_out_bits_4),
    .io_out_bits_5(memWriteDataMuxModule_io_out_bits_5),
    .io_out_bits_6(memWriteDataMuxModule_io_out_bits_6),
    .io_out_bits_7(memWriteDataMuxModule_io_out_bits_7),
    .io_out_bits_8(memWriteDataMuxModule_io_out_bits_8),
    .io_out_bits_9(memWriteDataMuxModule_io_out_bits_9),
    .io_out_bits_10(memWriteDataMuxModule_io_out_bits_10),
    .io_out_bits_11(memWriteDataMuxModule_io_out_bits_11),
    .io_out_bits_12(memWriteDataMuxModule_io_out_bits_12),
    .io_out_bits_13(memWriteDataMuxModule_io_out_bits_13),
    .io_out_bits_14(memWriteDataMuxModule_io_out_bits_14),
    .io_out_bits_15(memWriteDataMuxModule_io_out_bits_15),
    .io_out_bits_16(memWriteDataMuxModule_io_out_bits_16),
    .io_out_bits_17(memWriteDataMuxModule_io_out_bits_17),
    .io_out_bits_18(memWriteDataMuxModule_io_out_bits_18),
    .io_out_bits_19(memWriteDataMuxModule_io_out_bits_19),
    .io_out_bits_20(memWriteDataMuxModule_io_out_bits_20),
    .io_out_bits_21(memWriteDataMuxModule_io_out_bits_21),
    .io_out_bits_22(memWriteDataMuxModule_io_out_bits_22),
    .io_out_bits_23(memWriteDataMuxModule_io_out_bits_23),
    .io_out_bits_24(memWriteDataMuxModule_io_out_bits_24),
    .io_out_bits_25(memWriteDataMuxModule_io_out_bits_25),
    .io_out_bits_26(memWriteDataMuxModule_io_out_bits_26),
    .io_out_bits_27(memWriteDataMuxModule_io_out_bits_27),
    .io_out_bits_28(memWriteDataMuxModule_io_out_bits_28),
    .io_out_bits_29(memWriteDataMuxModule_io_out_bits_29),
    .io_out_bits_30(memWriteDataMuxModule_io_out_bits_30),
    .io_out_bits_31(memWriteDataMuxModule_io_out_bits_31)
  );
  Mux accWriteDataMuxModule ( // @[LocalRouter.scala 77:37]
    .io_in_0_ready(accWriteDataMuxModule_io_in_0_ready),
    .io_in_0_valid(accWriteDataMuxModule_io_in_0_valid),
    .io_in_0_bits_0(accWriteDataMuxModule_io_in_0_bits_0),
    .io_in_0_bits_1(accWriteDataMuxModule_io_in_0_bits_1),
    .io_in_0_bits_2(accWriteDataMuxModule_io_in_0_bits_2),
    .io_in_0_bits_3(accWriteDataMuxModule_io_in_0_bits_3),
    .io_in_0_bits_4(accWriteDataMuxModule_io_in_0_bits_4),
    .io_in_0_bits_5(accWriteDataMuxModule_io_in_0_bits_5),
    .io_in_0_bits_6(accWriteDataMuxModule_io_in_0_bits_6),
    .io_in_0_bits_7(accWriteDataMuxModule_io_in_0_bits_7),
    .io_in_0_bits_8(accWriteDataMuxModule_io_in_0_bits_8),
    .io_in_0_bits_9(accWriteDataMuxModule_io_in_0_bits_9),
    .io_in_0_bits_10(accWriteDataMuxModule_io_in_0_bits_10),
    .io_in_0_bits_11(accWriteDataMuxModule_io_in_0_bits_11),
    .io_in_0_bits_12(accWriteDataMuxModule_io_in_0_bits_12),
    .io_in_0_bits_13(accWriteDataMuxModule_io_in_0_bits_13),
    .io_in_0_bits_14(accWriteDataMuxModule_io_in_0_bits_14),
    .io_in_0_bits_15(accWriteDataMuxModule_io_in_0_bits_15),
    .io_in_0_bits_16(accWriteDataMuxModule_io_in_0_bits_16),
    .io_in_0_bits_17(accWriteDataMuxModule_io_in_0_bits_17),
    .io_in_0_bits_18(accWriteDataMuxModule_io_in_0_bits_18),
    .io_in_0_bits_19(accWriteDataMuxModule_io_in_0_bits_19),
    .io_in_0_bits_20(accWriteDataMuxModule_io_in_0_bits_20),
    .io_in_0_bits_21(accWriteDataMuxModule_io_in_0_bits_21),
    .io_in_0_bits_22(accWriteDataMuxModule_io_in_0_bits_22),
    .io_in_0_bits_23(accWriteDataMuxModule_io_in_0_bits_23),
    .io_in_0_bits_24(accWriteDataMuxModule_io_in_0_bits_24),
    .io_in_0_bits_25(accWriteDataMuxModule_io_in_0_bits_25),
    .io_in_0_bits_26(accWriteDataMuxModule_io_in_0_bits_26),
    .io_in_0_bits_27(accWriteDataMuxModule_io_in_0_bits_27),
    .io_in_0_bits_28(accWriteDataMuxModule_io_in_0_bits_28),
    .io_in_0_bits_29(accWriteDataMuxModule_io_in_0_bits_29),
    .io_in_0_bits_30(accWriteDataMuxModule_io_in_0_bits_30),
    .io_in_0_bits_31(accWriteDataMuxModule_io_in_0_bits_31),
    .io_in_1_ready(accWriteDataMuxModule_io_in_1_ready),
    .io_in_1_valid(accWriteDataMuxModule_io_in_1_valid),
    .io_in_1_bits_0(accWriteDataMuxModule_io_in_1_bits_0),
    .io_in_1_bits_1(accWriteDataMuxModule_io_in_1_bits_1),
    .io_in_1_bits_2(accWriteDataMuxModule_io_in_1_bits_2),
    .io_in_1_bits_3(accWriteDataMuxModule_io_in_1_bits_3),
    .io_in_1_bits_4(accWriteDataMuxModule_io_in_1_bits_4),
    .io_in_1_bits_5(accWriteDataMuxModule_io_in_1_bits_5),
    .io_in_1_bits_6(accWriteDataMuxModule_io_in_1_bits_6),
    .io_in_1_bits_7(accWriteDataMuxModule_io_in_1_bits_7),
    .io_in_1_bits_8(accWriteDataMuxModule_io_in_1_bits_8),
    .io_in_1_bits_9(accWriteDataMuxModule_io_in_1_bits_9),
    .io_in_1_bits_10(accWriteDataMuxModule_io_in_1_bits_10),
    .io_in_1_bits_11(accWriteDataMuxModule_io_in_1_bits_11),
    .io_in_1_bits_12(accWriteDataMuxModule_io_in_1_bits_12),
    .io_in_1_bits_13(accWriteDataMuxModule_io_in_1_bits_13),
    .io_in_1_bits_14(accWriteDataMuxModule_io_in_1_bits_14),
    .io_in_1_bits_15(accWriteDataMuxModule_io_in_1_bits_15),
    .io_in_1_bits_16(accWriteDataMuxModule_io_in_1_bits_16),
    .io_in_1_bits_17(accWriteDataMuxModule_io_in_1_bits_17),
    .io_in_1_bits_18(accWriteDataMuxModule_io_in_1_bits_18),
    .io_in_1_bits_19(accWriteDataMuxModule_io_in_1_bits_19),
    .io_in_1_bits_20(accWriteDataMuxModule_io_in_1_bits_20),
    .io_in_1_bits_21(accWriteDataMuxModule_io_in_1_bits_21),
    .io_in_1_bits_22(accWriteDataMuxModule_io_in_1_bits_22),
    .io_in_1_bits_23(accWriteDataMuxModule_io_in_1_bits_23),
    .io_in_1_bits_24(accWriteDataMuxModule_io_in_1_bits_24),
    .io_in_1_bits_25(accWriteDataMuxModule_io_in_1_bits_25),
    .io_in_1_bits_26(accWriteDataMuxModule_io_in_1_bits_26),
    .io_in_1_bits_27(accWriteDataMuxModule_io_in_1_bits_27),
    .io_in_1_bits_28(accWriteDataMuxModule_io_in_1_bits_28),
    .io_in_1_bits_29(accWriteDataMuxModule_io_in_1_bits_29),
    .io_in_1_bits_30(accWriteDataMuxModule_io_in_1_bits_30),
    .io_in_1_bits_31(accWriteDataMuxModule_io_in_1_bits_31),
    .io_sel_ready(accWriteDataMuxModule_io_sel_ready),
    .io_sel_valid(accWriteDataMuxModule_io_sel_valid),
    .io_sel_bits(accWriteDataMuxModule_io_sel_bits),
    .io_out_ready(accWriteDataMuxModule_io_out_ready),
    .io_out_valid(accWriteDataMuxModule_io_out_valid),
    .io_out_bits_0(accWriteDataMuxModule_io_out_bits_0),
    .io_out_bits_1(accWriteDataMuxModule_io_out_bits_1),
    .io_out_bits_2(accWriteDataMuxModule_io_out_bits_2),
    .io_out_bits_3(accWriteDataMuxModule_io_out_bits_3),
    .io_out_bits_4(accWriteDataMuxModule_io_out_bits_4),
    .io_out_bits_5(accWriteDataMuxModule_io_out_bits_5),
    .io_out_bits_6(accWriteDataMuxModule_io_out_bits_6),
    .io_out_bits_7(accWriteDataMuxModule_io_out_bits_7),
    .io_out_bits_8(accWriteDataMuxModule_io_out_bits_8),
    .io_out_bits_9(accWriteDataMuxModule_io_out_bits_9),
    .io_out_bits_10(accWriteDataMuxModule_io_out_bits_10),
    .io_out_bits_11(accWriteDataMuxModule_io_out_bits_11),
    .io_out_bits_12(accWriteDataMuxModule_io_out_bits_12),
    .io_out_bits_13(accWriteDataMuxModule_io_out_bits_13),
    .io_out_bits_14(accWriteDataMuxModule_io_out_bits_14),
    .io_out_bits_15(accWriteDataMuxModule_io_out_bits_15),
    .io_out_bits_16(accWriteDataMuxModule_io_out_bits_16),
    .io_out_bits_17(accWriteDataMuxModule_io_out_bits_17),
    .io_out_bits_18(accWriteDataMuxModule_io_out_bits_18),
    .io_out_bits_19(accWriteDataMuxModule_io_out_bits_19),
    .io_out_bits_20(accWriteDataMuxModule_io_out_bits_20),
    .io_out_bits_21(accWriteDataMuxModule_io_out_bits_21),
    .io_out_bits_22(accWriteDataMuxModule_io_out_bits_22),
    .io_out_bits_23(accWriteDataMuxModule_io_out_bits_23),
    .io_out_bits_24(accWriteDataMuxModule_io_out_bits_24),
    .io_out_bits_25(accWriteDataMuxModule_io_out_bits_25),
    .io_out_bits_26(accWriteDataMuxModule_io_out_bits_26),
    .io_out_bits_27(accWriteDataMuxModule_io_out_bits_27),
    .io_out_bits_28(accWriteDataMuxModule_io_out_bits_28),
    .io_out_bits_29(accWriteDataMuxModule_io_out_bits_29),
    .io_out_bits_30(accWriteDataMuxModule_io_out_bits_30),
    .io_out_bits_31(accWriteDataMuxModule_io_out_bits_31)
  );
  SizeHandler_2 sizeHandler ( // @[package.scala 33:29]
    .clock(sizeHandler_clock),
    .reset(sizeHandler_reset),
    .io_in_ready(sizeHandler_io_in_ready),
    .io_in_valid(sizeHandler_io_in_valid),
    .io_in_bits_sel(sizeHandler_io_in_bits_sel),
    .io_in_bits_size(sizeHandler_io_in_bits_size),
    .io_out_ready(sizeHandler_io_out_ready),
    .io_out_valid(sizeHandler_io_out_valid),
    .io_out_bits_sel(sizeHandler_io_out_bits_sel)
  );
  Queue_25 memReadDataDemux ( // @[Mem.scala 22:19]
    .clock(memReadDataDemux_clock),
    .reset(memReadDataDemux_reset),
    .io_enq_ready(memReadDataDemux_io_enq_ready),
    .io_enq_valid(memReadDataDemux_io_enq_valid),
    .io_enq_bits_sel(memReadDataDemux_io_enq_bits_sel),
    .io_enq_bits_size(memReadDataDemux_io_enq_bits_size),
    .io_deq_ready(memReadDataDemux_io_deq_ready),
    .io_deq_valid(memReadDataDemux_io_deq_valid),
    .io_deq_bits_sel(memReadDataDemux_io_deq_bits_sel),
    .io_deq_bits_size(memReadDataDemux_io_deq_bits_size)
  );
  SizeHandler_3 sizeHandler_1 ( // @[package.scala 33:29]
    .clock(sizeHandler_1_clock),
    .reset(sizeHandler_1_reset),
    .io_in_ready(sizeHandler_1_io_in_ready),
    .io_in_valid(sizeHandler_1_io_in_valid),
    .io_in_bits_sel(sizeHandler_1_io_in_bits_sel),
    .io_in_bits_size(sizeHandler_1_io_in_bits_size),
    .io_out_ready(sizeHandler_1_io_out_ready),
    .io_out_valid(sizeHandler_1_io_out_valid),
    .io_out_bits_sel(sizeHandler_1_io_out_bits_sel)
  );
  Queue_26 memWriteDataMux ( // @[Mem.scala 22:19]
    .clock(memWriteDataMux_clock),
    .reset(memWriteDataMux_reset),
    .io_enq_ready(memWriteDataMux_io_enq_ready),
    .io_enq_valid(memWriteDataMux_io_enq_valid),
    .io_enq_bits_sel(memWriteDataMux_io_enq_bits_sel),
    .io_enq_bits_size(memWriteDataMux_io_enq_bits_size),
    .io_deq_ready(memWriteDataMux_io_deq_ready),
    .io_deq_valid(memWriteDataMux_io_deq_valid),
    .io_deq_bits_sel(memWriteDataMux_io_deq_bits_sel),
    .io_deq_bits_size(memWriteDataMux_io_deq_bits_size)
  );
  SizeHandler_3 sizeHandler_2 ( // @[package.scala 33:29]
    .clock(sizeHandler_2_clock),
    .reset(sizeHandler_2_reset),
    .io_in_ready(sizeHandler_2_io_in_ready),
    .io_in_valid(sizeHandler_2_io_in_valid),
    .io_in_bits_sel(sizeHandler_2_io_in_bits_sel),
    .io_in_bits_size(sizeHandler_2_io_in_bits_size),
    .io_out_ready(sizeHandler_2_io_out_ready),
    .io_out_valid(sizeHandler_2_io_out_valid),
    .io_out_bits_sel(sizeHandler_2_io_out_bits_sel)
  );
  Queue_27 accWriteDataMux ( // @[Mem.scala 22:19]
    .clock(accWriteDataMux_clock),
    .reset(accWriteDataMux_reset),
    .io_enq_ready(accWriteDataMux_io_enq_ready),
    .io_enq_valid(accWriteDataMux_io_enq_valid),
    .io_enq_bits_sel(accWriteDataMux_io_enq_bits_sel),
    .io_enq_bits_size(accWriteDataMux_io_enq_bits_size),
    .io_deq_ready(accWriteDataMux_io_deq_ready),
    .io_deq_valid(accWriteDataMux_io_deq_valid),
    .io_deq_bits_sel(accWriteDataMux_io_deq_bits_sel),
    .io_deq_bits_size(accWriteDataMux_io_deq_bits_size)
  );
  MultiEnqueue enqueuer1 ( // @[MultiEnqueue.scala 182:43]
    .clock(enqueuer1_clock),
    .reset(enqueuer1_reset),
    .io_in_ready(enqueuer1_io_in_ready),
    .io_in_valid(enqueuer1_io_in_valid),
    .io_out_0_ready(enqueuer1_io_out_0_ready),
    .io_out_0_valid(enqueuer1_io_out_0_valid)
  );
  MultiEnqueue_1 enqueuer2 ( // @[MultiEnqueue.scala 182:43]
    .clock(enqueuer2_clock),
    .reset(enqueuer2_reset),
    .io_in_ready(enqueuer2_io_in_ready),
    .io_in_valid(enqueuer2_io_in_valid),
    .io_out_0_ready(enqueuer2_io_out_0_ready),
    .io_out_0_valid(enqueuer2_io_out_0_valid),
    .io_out_1_ready(enqueuer2_io_out_1_ready),
    .io_out_1_valid(enqueuer2_io_out_1_valid)
  );
  assign io_control_ready = io_control_bits_kind == 4'h1 ? enqueuer1_io_in_ready : _GEN_49; // @[LocalRouter.scala 123:72 124:19]
  assign io_mem_output_ready = memReadDataDemuxModule_io_in_ready; // @[LocalRouter.scala 62:32]
  assign io_mem_input_valid = memWriteDataMuxModule_io_out_valid; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_0 = memWriteDataMuxModule_io_out_bits_0; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_1 = memWriteDataMuxModule_io_out_bits_1; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_2 = memWriteDataMuxModule_io_out_bits_2; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_3 = memWriteDataMuxModule_io_out_bits_3; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_4 = memWriteDataMuxModule_io_out_bits_4; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_5 = memWriteDataMuxModule_io_out_bits_5; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_6 = memWriteDataMuxModule_io_out_bits_6; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_7 = memWriteDataMuxModule_io_out_bits_7; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_8 = memWriteDataMuxModule_io_out_bits_8; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_9 = memWriteDataMuxModule_io_out_bits_9; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_10 = memWriteDataMuxModule_io_out_bits_10; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_11 = memWriteDataMuxModule_io_out_bits_11; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_12 = memWriteDataMuxModule_io_out_bits_12; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_13 = memWriteDataMuxModule_io_out_bits_13; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_14 = memWriteDataMuxModule_io_out_bits_14; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_15 = memWriteDataMuxModule_io_out_bits_15; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_16 = memWriteDataMuxModule_io_out_bits_16; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_17 = memWriteDataMuxModule_io_out_bits_17; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_18 = memWriteDataMuxModule_io_out_bits_18; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_19 = memWriteDataMuxModule_io_out_bits_19; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_20 = memWriteDataMuxModule_io_out_bits_20; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_21 = memWriteDataMuxModule_io_out_bits_21; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_22 = memWriteDataMuxModule_io_out_bits_22; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_23 = memWriteDataMuxModule_io_out_bits_23; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_24 = memWriteDataMuxModule_io_out_bits_24; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_25 = memWriteDataMuxModule_io_out_bits_25; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_26 = memWriteDataMuxModule_io_out_bits_26; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_27 = memWriteDataMuxModule_io_out_bits_27; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_28 = memWriteDataMuxModule_io_out_bits_28; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_29 = memWriteDataMuxModule_io_out_bits_29; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_30 = memWriteDataMuxModule_io_out_bits_30; // @[LocalRouter.scala 75:16]
  assign io_mem_input_bits_31 = memWriteDataMuxModule_io_out_bits_31; // @[LocalRouter.scala 75:16]
  assign io_array_input_valid = memReadDataDemuxModule_io_out_1_valid; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_0 = memReadDataDemuxModule_io_out_1_bits_0; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_1 = memReadDataDemuxModule_io_out_1_bits_1; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_2 = memReadDataDemuxModule_io_out_1_bits_2; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_3 = memReadDataDemuxModule_io_out_1_bits_3; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_4 = memReadDataDemuxModule_io_out_1_bits_4; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_5 = memReadDataDemuxModule_io_out_1_bits_5; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_6 = memReadDataDemuxModule_io_out_1_bits_6; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_7 = memReadDataDemuxModule_io_out_1_bits_7; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_8 = memReadDataDemuxModule_io_out_1_bits_8; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_9 = memReadDataDemuxModule_io_out_1_bits_9; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_10 = memReadDataDemuxModule_io_out_1_bits_10; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_11 = memReadDataDemuxModule_io_out_1_bits_11; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_12 = memReadDataDemuxModule_io_out_1_bits_12; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_13 = memReadDataDemuxModule_io_out_1_bits_13; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_14 = memReadDataDemuxModule_io_out_1_bits_14; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_15 = memReadDataDemuxModule_io_out_1_bits_15; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_16 = memReadDataDemuxModule_io_out_1_bits_16; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_17 = memReadDataDemuxModule_io_out_1_bits_17; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_18 = memReadDataDemuxModule_io_out_1_bits_18; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_19 = memReadDataDemuxModule_io_out_1_bits_19; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_20 = memReadDataDemuxModule_io_out_1_bits_20; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_21 = memReadDataDemuxModule_io_out_1_bits_21; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_22 = memReadDataDemuxModule_io_out_1_bits_22; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_23 = memReadDataDemuxModule_io_out_1_bits_23; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_24 = memReadDataDemuxModule_io_out_1_bits_24; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_25 = memReadDataDemuxModule_io_out_1_bits_25; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_26 = memReadDataDemuxModule_io_out_1_bits_26; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_27 = memReadDataDemuxModule_io_out_1_bits_27; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_28 = memReadDataDemuxModule_io_out_1_bits_28; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_29 = memReadDataDemuxModule_io_out_1_bits_29; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_30 = memReadDataDemuxModule_io_out_1_bits_30; // @[LocalRouter.scala 64:18]
  assign io_array_input_bits_31 = memReadDataDemuxModule_io_out_1_bits_31; // @[LocalRouter.scala 64:18]
  assign io_array_output_ready = accWriteDataMuxModule_io_in_0_ready; // @[LocalRouter.scala 84:34]
  assign io_array_weightInput_valid = memReadDataDemuxModule_io_out_0_valid; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_0 = memReadDataDemuxModule_io_out_0_bits_0; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_1 = memReadDataDemuxModule_io_out_0_bits_1; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_2 = memReadDataDemuxModule_io_out_0_bits_2; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_3 = memReadDataDemuxModule_io_out_0_bits_3; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_4 = memReadDataDemuxModule_io_out_0_bits_4; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_5 = memReadDataDemuxModule_io_out_0_bits_5; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_6 = memReadDataDemuxModule_io_out_0_bits_6; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_7 = memReadDataDemuxModule_io_out_0_bits_7; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_8 = memReadDataDemuxModule_io_out_0_bits_8; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_9 = memReadDataDemuxModule_io_out_0_bits_9; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_10 = memReadDataDemuxModule_io_out_0_bits_10; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_11 = memReadDataDemuxModule_io_out_0_bits_11; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_12 = memReadDataDemuxModule_io_out_0_bits_12; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_13 = memReadDataDemuxModule_io_out_0_bits_13; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_14 = memReadDataDemuxModule_io_out_0_bits_14; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_15 = memReadDataDemuxModule_io_out_0_bits_15; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_16 = memReadDataDemuxModule_io_out_0_bits_16; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_17 = memReadDataDemuxModule_io_out_0_bits_17; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_18 = memReadDataDemuxModule_io_out_0_bits_18; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_19 = memReadDataDemuxModule_io_out_0_bits_19; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_20 = memReadDataDemuxModule_io_out_0_bits_20; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_21 = memReadDataDemuxModule_io_out_0_bits_21; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_22 = memReadDataDemuxModule_io_out_0_bits_22; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_23 = memReadDataDemuxModule_io_out_0_bits_23; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_24 = memReadDataDemuxModule_io_out_0_bits_24; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_25 = memReadDataDemuxModule_io_out_0_bits_25; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_26 = memReadDataDemuxModule_io_out_0_bits_26; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_27 = memReadDataDemuxModule_io_out_0_bits_27; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_28 = memReadDataDemuxModule_io_out_0_bits_28; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_29 = memReadDataDemuxModule_io_out_0_bits_29; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_30 = memReadDataDemuxModule_io_out_0_bits_30; // @[LocalRouter.scala 63:24]
  assign io_array_weightInput_bits_31 = memReadDataDemuxModule_io_out_0_bits_31; // @[LocalRouter.scala 63:24]
  assign io_acc_output_ready = memWriteDataMuxModule_io_in_1_ready; // @[LocalRouter.scala 74:34]
  assign io_acc_input_valid = accWriteDataMuxModule_io_out_valid; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_0 = accWriteDataMuxModule_io_out_bits_0; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_1 = accWriteDataMuxModule_io_out_bits_1; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_2 = accWriteDataMuxModule_io_out_bits_2; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_3 = accWriteDataMuxModule_io_out_bits_3; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_4 = accWriteDataMuxModule_io_out_bits_4; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_5 = accWriteDataMuxModule_io_out_bits_5; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_6 = accWriteDataMuxModule_io_out_bits_6; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_7 = accWriteDataMuxModule_io_out_bits_7; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_8 = accWriteDataMuxModule_io_out_bits_8; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_9 = accWriteDataMuxModule_io_out_bits_9; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_10 = accWriteDataMuxModule_io_out_bits_10; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_11 = accWriteDataMuxModule_io_out_bits_11; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_12 = accWriteDataMuxModule_io_out_bits_12; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_13 = accWriteDataMuxModule_io_out_bits_13; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_14 = accWriteDataMuxModule_io_out_bits_14; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_15 = accWriteDataMuxModule_io_out_bits_15; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_16 = accWriteDataMuxModule_io_out_bits_16; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_17 = accWriteDataMuxModule_io_out_bits_17; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_18 = accWriteDataMuxModule_io_out_bits_18; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_19 = accWriteDataMuxModule_io_out_bits_19; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_20 = accWriteDataMuxModule_io_out_bits_20; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_21 = accWriteDataMuxModule_io_out_bits_21; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_22 = accWriteDataMuxModule_io_out_bits_22; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_23 = accWriteDataMuxModule_io_out_bits_23; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_24 = accWriteDataMuxModule_io_out_bits_24; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_25 = accWriteDataMuxModule_io_out_bits_25; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_26 = accWriteDataMuxModule_io_out_bits_26; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_27 = accWriteDataMuxModule_io_out_bits_27; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_28 = accWriteDataMuxModule_io_out_bits_28; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_29 = accWriteDataMuxModule_io_out_bits_29; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_30 = accWriteDataMuxModule_io_out_bits_30; // @[LocalRouter.scala 86:16]
  assign io_acc_input_bits_31 = accWriteDataMuxModule_io_out_bits_31; // @[LocalRouter.scala 86:16]
  assign memReadDataDemuxModule_io_in_valid = io_mem_output_valid; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_0 = io_mem_output_bits_0; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_1 = io_mem_output_bits_1; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_2 = io_mem_output_bits_2; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_3 = io_mem_output_bits_3; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_4 = io_mem_output_bits_4; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_5 = io_mem_output_bits_5; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_6 = io_mem_output_bits_6; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_7 = io_mem_output_bits_7; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_8 = io_mem_output_bits_8; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_9 = io_mem_output_bits_9; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_10 = io_mem_output_bits_10; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_11 = io_mem_output_bits_11; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_12 = io_mem_output_bits_12; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_13 = io_mem_output_bits_13; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_14 = io_mem_output_bits_14; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_15 = io_mem_output_bits_15; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_16 = io_mem_output_bits_16; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_17 = io_mem_output_bits_17; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_18 = io_mem_output_bits_18; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_19 = io_mem_output_bits_19; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_20 = io_mem_output_bits_20; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_21 = io_mem_output_bits_21; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_22 = io_mem_output_bits_22; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_23 = io_mem_output_bits_23; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_24 = io_mem_output_bits_24; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_25 = io_mem_output_bits_25; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_26 = io_mem_output_bits_26; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_27 = io_mem_output_bits_27; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_28 = io_mem_output_bits_28; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_29 = io_mem_output_bits_29; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_30 = io_mem_output_bits_30; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_in_bits_31 = io_mem_output_bits_31; // @[LocalRouter.scala 62:32]
  assign memReadDataDemuxModule_io_sel_valid = sizeHandler_io_out_valid; // @[package.scala 39:18]
  assign memReadDataDemuxModule_io_sel_bits = sizeHandler_io_out_bits_sel; // @[package.scala 38:17]
  assign memReadDataDemuxModule_io_out_0_ready = io_array_weightInput_ready; // @[LocalRouter.scala 63:24]
  assign memReadDataDemuxModule_io_out_1_ready = io_array_input_ready; // @[LocalRouter.scala 64:18]
  assign memReadDataDemuxModule_io_out_2_ready = accWriteDataMuxModule_io_in_1_ready; // @[LocalRouter.scala 85:34]
  assign memWriteDataMuxModule_io_in_0_valid = 1'h0; // @[package.scala 405:15]
  assign memWriteDataMuxModule_io_in_0_bits_0 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_1 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_2 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_3 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_4 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_5 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_6 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_7 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_8 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_9 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_10 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_11 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_12 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_13 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_14 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_15 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_16 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_17 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_18 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_19 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_20 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_21 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_22 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_23 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_24 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_25 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_26 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_27 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_28 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_29 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_30 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_0_bits_31 = 16'sh0; // @[package.scala 75:57]
  assign memWriteDataMuxModule_io_in_1_valid = io_acc_output_valid; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_0 = io_acc_output_bits_0; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_1 = io_acc_output_bits_1; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_2 = io_acc_output_bits_2; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_3 = io_acc_output_bits_3; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_4 = io_acc_output_bits_4; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_5 = io_acc_output_bits_5; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_6 = io_acc_output_bits_6; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_7 = io_acc_output_bits_7; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_8 = io_acc_output_bits_8; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_9 = io_acc_output_bits_9; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_10 = io_acc_output_bits_10; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_11 = io_acc_output_bits_11; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_12 = io_acc_output_bits_12; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_13 = io_acc_output_bits_13; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_14 = io_acc_output_bits_14; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_15 = io_acc_output_bits_15; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_16 = io_acc_output_bits_16; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_17 = io_acc_output_bits_17; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_18 = io_acc_output_bits_18; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_19 = io_acc_output_bits_19; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_20 = io_acc_output_bits_20; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_21 = io_acc_output_bits_21; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_22 = io_acc_output_bits_22; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_23 = io_acc_output_bits_23; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_24 = io_acc_output_bits_24; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_25 = io_acc_output_bits_25; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_26 = io_acc_output_bits_26; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_27 = io_acc_output_bits_27; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_28 = io_acc_output_bits_28; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_29 = io_acc_output_bits_29; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_30 = io_acc_output_bits_30; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_in_1_bits_31 = io_acc_output_bits_31; // @[LocalRouter.scala 74:34]
  assign memWriteDataMuxModule_io_sel_valid = sizeHandler_1_io_out_valid; // @[package.scala 39:18]
  assign memWriteDataMuxModule_io_sel_bits = sizeHandler_1_io_out_bits_sel; // @[package.scala 38:17]
  assign memWriteDataMuxModule_io_out_ready = io_mem_input_ready; // @[LocalRouter.scala 75:16]
  assign accWriteDataMuxModule_io_in_0_valid = io_array_output_valid; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_0 = io_array_output_bits_0; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_1 = io_array_output_bits_1; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_2 = io_array_output_bits_2; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_3 = io_array_output_bits_3; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_4 = io_array_output_bits_4; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_5 = io_array_output_bits_5; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_6 = io_array_output_bits_6; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_7 = io_array_output_bits_7; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_8 = io_array_output_bits_8; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_9 = io_array_output_bits_9; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_10 = io_array_output_bits_10; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_11 = io_array_output_bits_11; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_12 = io_array_output_bits_12; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_13 = io_array_output_bits_13; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_14 = io_array_output_bits_14; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_15 = io_array_output_bits_15; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_16 = io_array_output_bits_16; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_17 = io_array_output_bits_17; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_18 = io_array_output_bits_18; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_19 = io_array_output_bits_19; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_20 = io_array_output_bits_20; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_21 = io_array_output_bits_21; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_22 = io_array_output_bits_22; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_23 = io_array_output_bits_23; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_24 = io_array_output_bits_24; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_25 = io_array_output_bits_25; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_26 = io_array_output_bits_26; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_27 = io_array_output_bits_27; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_28 = io_array_output_bits_28; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_29 = io_array_output_bits_29; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_30 = io_array_output_bits_30; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_0_bits_31 = io_array_output_bits_31; // @[LocalRouter.scala 84:34]
  assign accWriteDataMuxModule_io_in_1_valid = memReadDataDemuxModule_io_out_2_valid; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_0 = memReadDataDemuxModule_io_out_2_bits_0; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_1 = memReadDataDemuxModule_io_out_2_bits_1; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_2 = memReadDataDemuxModule_io_out_2_bits_2; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_3 = memReadDataDemuxModule_io_out_2_bits_3; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_4 = memReadDataDemuxModule_io_out_2_bits_4; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_5 = memReadDataDemuxModule_io_out_2_bits_5; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_6 = memReadDataDemuxModule_io_out_2_bits_6; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_7 = memReadDataDemuxModule_io_out_2_bits_7; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_8 = memReadDataDemuxModule_io_out_2_bits_8; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_9 = memReadDataDemuxModule_io_out_2_bits_9; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_10 = memReadDataDemuxModule_io_out_2_bits_10; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_11 = memReadDataDemuxModule_io_out_2_bits_11; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_12 = memReadDataDemuxModule_io_out_2_bits_12; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_13 = memReadDataDemuxModule_io_out_2_bits_13; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_14 = memReadDataDemuxModule_io_out_2_bits_14; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_15 = memReadDataDemuxModule_io_out_2_bits_15; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_16 = memReadDataDemuxModule_io_out_2_bits_16; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_17 = memReadDataDemuxModule_io_out_2_bits_17; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_18 = memReadDataDemuxModule_io_out_2_bits_18; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_19 = memReadDataDemuxModule_io_out_2_bits_19; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_20 = memReadDataDemuxModule_io_out_2_bits_20; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_21 = memReadDataDemuxModule_io_out_2_bits_21; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_22 = memReadDataDemuxModule_io_out_2_bits_22; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_23 = memReadDataDemuxModule_io_out_2_bits_23; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_24 = memReadDataDemuxModule_io_out_2_bits_24; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_25 = memReadDataDemuxModule_io_out_2_bits_25; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_26 = memReadDataDemuxModule_io_out_2_bits_26; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_27 = memReadDataDemuxModule_io_out_2_bits_27; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_28 = memReadDataDemuxModule_io_out_2_bits_28; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_29 = memReadDataDemuxModule_io_out_2_bits_29; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_30 = memReadDataDemuxModule_io_out_2_bits_30; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_in_1_bits_31 = memReadDataDemuxModule_io_out_2_bits_31; // @[LocalRouter.scala 85:34]
  assign accWriteDataMuxModule_io_sel_valid = sizeHandler_2_io_out_valid; // @[package.scala 39:18]
  assign accWriteDataMuxModule_io_sel_bits = sizeHandler_2_io_out_bits_sel; // @[package.scala 38:17]
  assign accWriteDataMuxModule_io_out_ready = io_acc_input_ready; // @[LocalRouter.scala 86:16]
  assign sizeHandler_clock = clock;
  assign sizeHandler_reset = reset;
  assign sizeHandler_io_in_valid = memReadDataDemux_io_deq_valid; // @[Mem.scala 23:7]
  assign sizeHandler_io_in_bits_sel = memReadDataDemux_io_deq_bits_sel; // @[Mem.scala 23:7]
  assign sizeHandler_io_in_bits_size = memReadDataDemux_io_deq_bits_size; // @[Mem.scala 23:7]
  assign sizeHandler_io_out_ready = memReadDataDemuxModule_io_sel_ready; // @[package.scala 40:30]
  assign memReadDataDemux_clock = clock;
  assign memReadDataDemux_reset = reset;
  assign memReadDataDemux_io_enq_valid = io_control_bits_kind == 4'h1 ? io_control_ready_memWriteDataMux_io_enq_w_valid
     : _GEN_42; // @[LocalRouter.scala 123:72 MultiEnqueue.scala 61:10]
  assign memReadDataDemux_io_enq_bits_sel = io_control_bits_kind == 4'h1 ? 2'h0 : _GEN_43; // @[LocalRouter.scala 123:72 MultiEnqueue.scala 61:10]
  assign memReadDataDemux_io_enq_bits_size = io_control_bits_kind == 4'h1 ? io_control_bits_size : _GEN_44; // @[LocalRouter.scala 123:72 MultiEnqueue.scala 61:10]
  assign memReadDataDemux_io_deq_ready = sizeHandler_io_in_ready; // @[Mem.scala 23:7]
  assign sizeHandler_1_clock = clock;
  assign sizeHandler_1_reset = reset;
  assign sizeHandler_1_io_in_valid = memWriteDataMux_io_deq_valid; // @[Mem.scala 23:7]
  assign sizeHandler_1_io_in_bits_sel = memWriteDataMux_io_deq_bits_sel; // @[Mem.scala 23:7]
  assign sizeHandler_1_io_in_bits_size = memWriteDataMux_io_deq_bits_size; // @[Mem.scala 23:7]
  assign sizeHandler_1_io_out_ready = memWriteDataMuxModule_io_sel_ready; // @[package.scala 40:30]
  assign memWriteDataMux_clock = clock;
  assign memWriteDataMux_reset = reset;
  assign memWriteDataMux_io_enq_valid = io_control_bits_kind == 4'h1 ? 1'h0 : _GEN_52; // @[LocalRouter.scala 123:72 package.scala 405:15]
  assign memWriteDataMux_io_enq_bits_sel = io_control_bits_kind == 4'h1 ? 1'h0 : _GEN_53; // @[LocalRouter.scala 123:72 package.scala 404:14]
  assign memWriteDataMux_io_enq_bits_size = io_control_bits_kind == 4'h1 ? 14'h0 : _GEN_54; // @[LocalRouter.scala 123:72 package.scala 404:14]
  assign memWriteDataMux_io_deq_ready = sizeHandler_1_io_in_ready; // @[Mem.scala 23:7]
  assign sizeHandler_2_clock = clock;
  assign sizeHandler_2_reset = reset;
  assign sizeHandler_2_io_in_valid = accWriteDataMux_io_deq_valid; // @[Mem.scala 23:7]
  assign sizeHandler_2_io_in_bits_sel = accWriteDataMux_io_deq_bits_sel; // @[Mem.scala 23:7]
  assign sizeHandler_2_io_in_bits_size = accWriteDataMux_io_deq_bits_size; // @[Mem.scala 23:7]
  assign sizeHandler_2_io_out_ready = accWriteDataMuxModule_io_sel_ready; // @[package.scala 40:30]
  assign accWriteDataMux_clock = clock;
  assign accWriteDataMux_reset = reset;
  assign accWriteDataMux_io_enq_valid = io_control_bits_kind == 4'h1 ? 1'h0 : _GEN_46; // @[LocalRouter.scala 123:72 package.scala 405:15]
  assign accWriteDataMux_io_enq_bits_sel = io_control_bits_kind == 4'h1 ? 1'h0 : _GEN_47; // @[LocalRouter.scala 123:72 package.scala 404:14]
  assign accWriteDataMux_io_enq_bits_size = io_control_bits_kind == 4'h1 ? 14'h0 : _GEN_48; // @[LocalRouter.scala 123:72 package.scala 404:14]
  assign accWriteDataMux_io_deq_ready = sizeHandler_2_io_in_ready; // @[Mem.scala 23:7]
  assign enqueuer1_clock = clock;
  assign enqueuer1_reset = reset;
  assign enqueuer1_io_in_valid = io_control_bits_kind == 4'h1 ? io_control_valid : _GEN_50; // @[LocalRouter.scala 123:72 MultiEnqueue.scala 60:17]
  assign enqueuer1_io_out_0_ready = io_control_bits_kind == 4'h1 ? io_control_ready_memReadDataDemux_io_enq_w_2_ready :
    _GEN_51; // @[LocalRouter.scala 123:72 ReadyValid.scala 19:11]
  assign enqueuer2_clock = clock;
  assign enqueuer2_reset = reset;
  assign enqueuer2_io_in_valid = io_control_bits_kind == 4'h1 ? 1'h0 : _GEN_40; // @[LocalRouter.scala 123:72 MultiEnqueue.scala 40:17]
  assign enqueuer2_io_out_0_ready = io_control_bits_kind == 4'h1 ? 1'h0 : _GEN_41; // @[LocalRouter.scala 123:72 MultiEnqueue.scala 42:18]
  assign enqueuer2_io_out_1_ready = io_control_bits_kind == 4'h1 ? 1'h0 : _GEN_45; // @[LocalRouter.scala 123:72 MultiEnqueue.scala 42:18]
endmodule
module HostRouter(
  output        io_control_ready,
  input         io_control_valid,
  input  [1:0]  io_control_bits_kind,
  output        io_dram0_dataIn_ready,
  input         io_dram0_dataIn_valid,
  input  [15:0] io_dram0_dataIn_bits_0,
  input  [15:0] io_dram0_dataIn_bits_1,
  input  [15:0] io_dram0_dataIn_bits_2,
  input  [15:0] io_dram0_dataIn_bits_3,
  input  [15:0] io_dram0_dataIn_bits_4,
  input  [15:0] io_dram0_dataIn_bits_5,
  input  [15:0] io_dram0_dataIn_bits_6,
  input  [15:0] io_dram0_dataIn_bits_7,
  input  [15:0] io_dram0_dataIn_bits_8,
  input  [15:0] io_dram0_dataIn_bits_9,
  input  [15:0] io_dram0_dataIn_bits_10,
  input  [15:0] io_dram0_dataIn_bits_11,
  input  [15:0] io_dram0_dataIn_bits_12,
  input  [15:0] io_dram0_dataIn_bits_13,
  input  [15:0] io_dram0_dataIn_bits_14,
  input  [15:0] io_dram0_dataIn_bits_15,
  input  [15:0] io_dram0_dataIn_bits_16,
  input  [15:0] io_dram0_dataIn_bits_17,
  input  [15:0] io_dram0_dataIn_bits_18,
  input  [15:0] io_dram0_dataIn_bits_19,
  input  [15:0] io_dram0_dataIn_bits_20,
  input  [15:0] io_dram0_dataIn_bits_21,
  input  [15:0] io_dram0_dataIn_bits_22,
  input  [15:0] io_dram0_dataIn_bits_23,
  input  [15:0] io_dram0_dataIn_bits_24,
  input  [15:0] io_dram0_dataIn_bits_25,
  input  [15:0] io_dram0_dataIn_bits_26,
  input  [15:0] io_dram0_dataIn_bits_27,
  input  [15:0] io_dram0_dataIn_bits_28,
  input  [15:0] io_dram0_dataIn_bits_29,
  input  [15:0] io_dram0_dataIn_bits_30,
  input  [15:0] io_dram0_dataIn_bits_31,
  input         io_dram0_dataOut_ready,
  output        io_dram0_dataOut_valid,
  output [15:0] io_dram0_dataOut_bits_0,
  output [15:0] io_dram0_dataOut_bits_1,
  output [15:0] io_dram0_dataOut_bits_2,
  output [15:0] io_dram0_dataOut_bits_3,
  output [15:0] io_dram0_dataOut_bits_4,
  output [15:0] io_dram0_dataOut_bits_5,
  output [15:0] io_dram0_dataOut_bits_6,
  output [15:0] io_dram0_dataOut_bits_7,
  output [15:0] io_dram0_dataOut_bits_8,
  output [15:0] io_dram0_dataOut_bits_9,
  output [15:0] io_dram0_dataOut_bits_10,
  output [15:0] io_dram0_dataOut_bits_11,
  output [15:0] io_dram0_dataOut_bits_12,
  output [15:0] io_dram0_dataOut_bits_13,
  output [15:0] io_dram0_dataOut_bits_14,
  output [15:0] io_dram0_dataOut_bits_15,
  output [15:0] io_dram0_dataOut_bits_16,
  output [15:0] io_dram0_dataOut_bits_17,
  output [15:0] io_dram0_dataOut_bits_18,
  output [15:0] io_dram0_dataOut_bits_19,
  output [15:0] io_dram0_dataOut_bits_20,
  output [15:0] io_dram0_dataOut_bits_21,
  output [15:0] io_dram0_dataOut_bits_22,
  output [15:0] io_dram0_dataOut_bits_23,
  output [15:0] io_dram0_dataOut_bits_24,
  output [15:0] io_dram0_dataOut_bits_25,
  output [15:0] io_dram0_dataOut_bits_26,
  output [15:0] io_dram0_dataOut_bits_27,
  output [15:0] io_dram0_dataOut_bits_28,
  output [15:0] io_dram0_dataOut_bits_29,
  output [15:0] io_dram0_dataOut_bits_30,
  output [15:0] io_dram0_dataOut_bits_31,
  output        io_dram1_dataIn_ready,
  input         io_dram1_dataIn_valid,
  input  [15:0] io_dram1_dataIn_bits_0,
  input  [15:0] io_dram1_dataIn_bits_1,
  input  [15:0] io_dram1_dataIn_bits_2,
  input  [15:0] io_dram1_dataIn_bits_3,
  input  [15:0] io_dram1_dataIn_bits_4,
  input  [15:0] io_dram1_dataIn_bits_5,
  input  [15:0] io_dram1_dataIn_bits_6,
  input  [15:0] io_dram1_dataIn_bits_7,
  input  [15:0] io_dram1_dataIn_bits_8,
  input  [15:0] io_dram1_dataIn_bits_9,
  input  [15:0] io_dram1_dataIn_bits_10,
  input  [15:0] io_dram1_dataIn_bits_11,
  input  [15:0] io_dram1_dataIn_bits_12,
  input  [15:0] io_dram1_dataIn_bits_13,
  input  [15:0] io_dram1_dataIn_bits_14,
  input  [15:0] io_dram1_dataIn_bits_15,
  input  [15:0] io_dram1_dataIn_bits_16,
  input  [15:0] io_dram1_dataIn_bits_17,
  input  [15:0] io_dram1_dataIn_bits_18,
  input  [15:0] io_dram1_dataIn_bits_19,
  input  [15:0] io_dram1_dataIn_bits_20,
  input  [15:0] io_dram1_dataIn_bits_21,
  input  [15:0] io_dram1_dataIn_bits_22,
  input  [15:0] io_dram1_dataIn_bits_23,
  input  [15:0] io_dram1_dataIn_bits_24,
  input  [15:0] io_dram1_dataIn_bits_25,
  input  [15:0] io_dram1_dataIn_bits_26,
  input  [15:0] io_dram1_dataIn_bits_27,
  input  [15:0] io_dram1_dataIn_bits_28,
  input  [15:0] io_dram1_dataIn_bits_29,
  input  [15:0] io_dram1_dataIn_bits_30,
  input  [15:0] io_dram1_dataIn_bits_31,
  input         io_dram1_dataOut_ready,
  output        io_dram1_dataOut_valid,
  output [15:0] io_dram1_dataOut_bits_0,
  output [15:0] io_dram1_dataOut_bits_1,
  output [15:0] io_dram1_dataOut_bits_2,
  output [15:0] io_dram1_dataOut_bits_3,
  output [15:0] io_dram1_dataOut_bits_4,
  output [15:0] io_dram1_dataOut_bits_5,
  output [15:0] io_dram1_dataOut_bits_6,
  output [15:0] io_dram1_dataOut_bits_7,
  output [15:0] io_dram1_dataOut_bits_8,
  output [15:0] io_dram1_dataOut_bits_9,
  output [15:0] io_dram1_dataOut_bits_10,
  output [15:0] io_dram1_dataOut_bits_11,
  output [15:0] io_dram1_dataOut_bits_12,
  output [15:0] io_dram1_dataOut_bits_13,
  output [15:0] io_dram1_dataOut_bits_14,
  output [15:0] io_dram1_dataOut_bits_15,
  output [15:0] io_dram1_dataOut_bits_16,
  output [15:0] io_dram1_dataOut_bits_17,
  output [15:0] io_dram1_dataOut_bits_18,
  output [15:0] io_dram1_dataOut_bits_19,
  output [15:0] io_dram1_dataOut_bits_20,
  output [15:0] io_dram1_dataOut_bits_21,
  output [15:0] io_dram1_dataOut_bits_22,
  output [15:0] io_dram1_dataOut_bits_23,
  output [15:0] io_dram1_dataOut_bits_24,
  output [15:0] io_dram1_dataOut_bits_25,
  output [15:0] io_dram1_dataOut_bits_26,
  output [15:0] io_dram1_dataOut_bits_27,
  output [15:0] io_dram1_dataOut_bits_28,
  output [15:0] io_dram1_dataOut_bits_29,
  output [15:0] io_dram1_dataOut_bits_30,
  output [15:0] io_dram1_dataOut_bits_31,
  output        io_mem_output_ready,
  input         io_mem_output_valid,
  input  [15:0] io_mem_output_bits_0,
  input  [15:0] io_mem_output_bits_1,
  input  [15:0] io_mem_output_bits_2,
  input  [15:0] io_mem_output_bits_3,
  input  [15:0] io_mem_output_bits_4,
  input  [15:0] io_mem_output_bits_5,
  input  [15:0] io_mem_output_bits_6,
  input  [15:0] io_mem_output_bits_7,
  input  [15:0] io_mem_output_bits_8,
  input  [15:0] io_mem_output_bits_9,
  input  [15:0] io_mem_output_bits_10,
  input  [15:0] io_mem_output_bits_11,
  input  [15:0] io_mem_output_bits_12,
  input  [15:0] io_mem_output_bits_13,
  input  [15:0] io_mem_output_bits_14,
  input  [15:0] io_mem_output_bits_15,
  input  [15:0] io_mem_output_bits_16,
  input  [15:0] io_mem_output_bits_17,
  input  [15:0] io_mem_output_bits_18,
  input  [15:0] io_mem_output_bits_19,
  input  [15:0] io_mem_output_bits_20,
  input  [15:0] io_mem_output_bits_21,
  input  [15:0] io_mem_output_bits_22,
  input  [15:0] io_mem_output_bits_23,
  input  [15:0] io_mem_output_bits_24,
  input  [15:0] io_mem_output_bits_25,
  input  [15:0] io_mem_output_bits_26,
  input  [15:0] io_mem_output_bits_27,
  input  [15:0] io_mem_output_bits_28,
  input  [15:0] io_mem_output_bits_29,
  input  [15:0] io_mem_output_bits_30,
  input  [15:0] io_mem_output_bits_31,
  input         io_mem_input_ready,
  output        io_mem_input_valid,
  output [15:0] io_mem_input_bits_0,
  output [15:0] io_mem_input_bits_1,
  output [15:0] io_mem_input_bits_2,
  output [15:0] io_mem_input_bits_3,
  output [15:0] io_mem_input_bits_4,
  output [15:0] io_mem_input_bits_5,
  output [15:0] io_mem_input_bits_6,
  output [15:0] io_mem_input_bits_7,
  output [15:0] io_mem_input_bits_8,
  output [15:0] io_mem_input_bits_9,
  output [15:0] io_mem_input_bits_10,
  output [15:0] io_mem_input_bits_11,
  output [15:0] io_mem_input_bits_12,
  output [15:0] io_mem_input_bits_13,
  output [15:0] io_mem_input_bits_14,
  output [15:0] io_mem_input_bits_15,
  output [15:0] io_mem_input_bits_16,
  output [15:0] io_mem_input_bits_17,
  output [15:0] io_mem_input_bits_18,
  output [15:0] io_mem_input_bits_19,
  output [15:0] io_mem_input_bits_20,
  output [15:0] io_mem_input_bits_21,
  output [15:0] io_mem_input_bits_22,
  output [15:0] io_mem_input_bits_23,
  output [15:0] io_mem_input_bits_24,
  output [15:0] io_mem_input_bits_25,
  output [15:0] io_mem_input_bits_26,
  output [15:0] io_mem_input_bits_27,
  output [15:0] io_mem_input_bits_28,
  output [15:0] io_mem_input_bits_29,
  output [15:0] io_mem_input_bits_30,
  output [15:0] io_mem_input_bits_31
);
  wire  dataIn_mux_io_in_0_ready; // @[Mux.scala 71:21]
  wire  dataIn_mux_io_in_0_valid; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_0; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_1; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_2; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_3; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_4; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_5; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_6; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_7; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_8; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_9; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_10; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_11; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_12; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_13; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_14; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_15; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_16; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_17; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_18; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_19; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_20; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_21; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_22; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_23; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_24; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_25; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_26; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_27; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_28; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_29; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_30; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_0_bits_31; // @[Mux.scala 71:21]
  wire  dataIn_mux_io_in_1_ready; // @[Mux.scala 71:21]
  wire  dataIn_mux_io_in_1_valid; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_0; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_1; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_2; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_3; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_4; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_5; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_6; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_7; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_8; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_9; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_10; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_11; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_12; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_13; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_14; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_15; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_16; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_17; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_18; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_19; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_20; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_21; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_22; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_23; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_24; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_25; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_26; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_27; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_28; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_29; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_30; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_in_1_bits_31; // @[Mux.scala 71:21]
  wire  dataIn_mux_io_sel_ready; // @[Mux.scala 71:21]
  wire  dataIn_mux_io_sel_valid; // @[Mux.scala 71:21]
  wire  dataIn_mux_io_sel_bits; // @[Mux.scala 71:21]
  wire  dataIn_mux_io_out_ready; // @[Mux.scala 71:21]
  wire  dataIn_mux_io_out_valid; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_0; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_1; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_2; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_3; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_4; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_5; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_6; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_7; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_8; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_9; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_10; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_11; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_12; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_13; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_14; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_15; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_16; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_17; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_18; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_19; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_20; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_21; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_22; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_23; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_24; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_25; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_26; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_27; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_28; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_29; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_30; // @[Mux.scala 71:21]
  wire [15:0] dataIn_mux_io_out_bits_31; // @[Mux.scala 71:21]
  wire  dataOut_demux_io_in_ready; // @[Demux.scala 46:23]
  wire  dataOut_demux_io_in_valid; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_0; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_1; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_2; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_3; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_4; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_5; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_6; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_7; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_8; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_9; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_10; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_11; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_12; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_13; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_14; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_15; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_16; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_17; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_18; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_19; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_20; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_21; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_22; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_23; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_24; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_25; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_26; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_27; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_28; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_29; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_30; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_in_bits_31; // @[Demux.scala 46:23]
  wire  dataOut_demux_io_sel_ready; // @[Demux.scala 46:23]
  wire  dataOut_demux_io_sel_valid; // @[Demux.scala 46:23]
  wire  dataOut_demux_io_sel_bits; // @[Demux.scala 46:23]
  wire  dataOut_demux_io_out_0_ready; // @[Demux.scala 46:23]
  wire  dataOut_demux_io_out_0_valid; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_0; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_1; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_2; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_3; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_4; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_5; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_6; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_7; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_8; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_9; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_10; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_11; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_12; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_13; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_14; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_15; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_16; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_17; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_18; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_19; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_20; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_21; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_22; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_23; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_24; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_25; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_26; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_27; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_28; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_29; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_30; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_0_bits_31; // @[Demux.scala 46:23]
  wire  dataOut_demux_io_out_1_ready; // @[Demux.scala 46:23]
  wire  dataOut_demux_io_out_1_valid; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_0; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_1; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_2; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_3; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_4; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_5; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_6; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_7; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_8; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_9; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_10; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_11; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_12; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_13; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_14; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_15; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_16; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_17; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_18; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_19; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_20; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_21; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_22; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_23; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_24; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_25; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_26; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_27; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_28; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_29; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_30; // @[Demux.scala 46:23]
  wire [15:0] dataOut_demux_io_out_1_bits_31; // @[Demux.scala 46:23]
  wire  isDataIn = io_control_bits_kind == 2'h0 | io_control_bits_kind == 2'h2; // @[HostRouter.scala 57:18]
  wire  isDataOut = io_control_bits_kind == 2'h1 | io_control_bits_kind == 2'h3; // @[HostRouter.scala 61:19]
  Mux dataIn_mux ( // @[Mux.scala 71:21]
    .io_in_0_ready(dataIn_mux_io_in_0_ready),
    .io_in_0_valid(dataIn_mux_io_in_0_valid),
    .io_in_0_bits_0(dataIn_mux_io_in_0_bits_0),
    .io_in_0_bits_1(dataIn_mux_io_in_0_bits_1),
    .io_in_0_bits_2(dataIn_mux_io_in_0_bits_2),
    .io_in_0_bits_3(dataIn_mux_io_in_0_bits_3),
    .io_in_0_bits_4(dataIn_mux_io_in_0_bits_4),
    .io_in_0_bits_5(dataIn_mux_io_in_0_bits_5),
    .io_in_0_bits_6(dataIn_mux_io_in_0_bits_6),
    .io_in_0_bits_7(dataIn_mux_io_in_0_bits_7),
    .io_in_0_bits_8(dataIn_mux_io_in_0_bits_8),
    .io_in_0_bits_9(dataIn_mux_io_in_0_bits_9),
    .io_in_0_bits_10(dataIn_mux_io_in_0_bits_10),
    .io_in_0_bits_11(dataIn_mux_io_in_0_bits_11),
    .io_in_0_bits_12(dataIn_mux_io_in_0_bits_12),
    .io_in_0_bits_13(dataIn_mux_io_in_0_bits_13),
    .io_in_0_bits_14(dataIn_mux_io_in_0_bits_14),
    .io_in_0_bits_15(dataIn_mux_io_in_0_bits_15),
    .io_in_0_bits_16(dataIn_mux_io_in_0_bits_16),
    .io_in_0_bits_17(dataIn_mux_io_in_0_bits_17),
    .io_in_0_bits_18(dataIn_mux_io_in_0_bits_18),
    .io_in_0_bits_19(dataIn_mux_io_in_0_bits_19),
    .io_in_0_bits_20(dataIn_mux_io_in_0_bits_20),
    .io_in_0_bits_21(dataIn_mux_io_in_0_bits_21),
    .io_in_0_bits_22(dataIn_mux_io_in_0_bits_22),
    .io_in_0_bits_23(dataIn_mux_io_in_0_bits_23),
    .io_in_0_bits_24(dataIn_mux_io_in_0_bits_24),
    .io_in_0_bits_25(dataIn_mux_io_in_0_bits_25),
    .io_in_0_bits_26(dataIn_mux_io_in_0_bits_26),
    .io_in_0_bits_27(dataIn_mux_io_in_0_bits_27),
    .io_in_0_bits_28(dataIn_mux_io_in_0_bits_28),
    .io_in_0_bits_29(dataIn_mux_io_in_0_bits_29),
    .io_in_0_bits_30(dataIn_mux_io_in_0_bits_30),
    .io_in_0_bits_31(dataIn_mux_io_in_0_bits_31),
    .io_in_1_ready(dataIn_mux_io_in_1_ready),
    .io_in_1_valid(dataIn_mux_io_in_1_valid),
    .io_in_1_bits_0(dataIn_mux_io_in_1_bits_0),
    .io_in_1_bits_1(dataIn_mux_io_in_1_bits_1),
    .io_in_1_bits_2(dataIn_mux_io_in_1_bits_2),
    .io_in_1_bits_3(dataIn_mux_io_in_1_bits_3),
    .io_in_1_bits_4(dataIn_mux_io_in_1_bits_4),
    .io_in_1_bits_5(dataIn_mux_io_in_1_bits_5),
    .io_in_1_bits_6(dataIn_mux_io_in_1_bits_6),
    .io_in_1_bits_7(dataIn_mux_io_in_1_bits_7),
    .io_in_1_bits_8(dataIn_mux_io_in_1_bits_8),
    .io_in_1_bits_9(dataIn_mux_io_in_1_bits_9),
    .io_in_1_bits_10(dataIn_mux_io_in_1_bits_10),
    .io_in_1_bits_11(dataIn_mux_io_in_1_bits_11),
    .io_in_1_bits_12(dataIn_mux_io_in_1_bits_12),
    .io_in_1_bits_13(dataIn_mux_io_in_1_bits_13),
    .io_in_1_bits_14(dataIn_mux_io_in_1_bits_14),
    .io_in_1_bits_15(dataIn_mux_io_in_1_bits_15),
    .io_in_1_bits_16(dataIn_mux_io_in_1_bits_16),
    .io_in_1_bits_17(dataIn_mux_io_in_1_bits_17),
    .io_in_1_bits_18(dataIn_mux_io_in_1_bits_18),
    .io_in_1_bits_19(dataIn_mux_io_in_1_bits_19),
    .io_in_1_bits_20(dataIn_mux_io_in_1_bits_20),
    .io_in_1_bits_21(dataIn_mux_io_in_1_bits_21),
    .io_in_1_bits_22(dataIn_mux_io_in_1_bits_22),
    .io_in_1_bits_23(dataIn_mux_io_in_1_bits_23),
    .io_in_1_bits_24(dataIn_mux_io_in_1_bits_24),
    .io_in_1_bits_25(dataIn_mux_io_in_1_bits_25),
    .io_in_1_bits_26(dataIn_mux_io_in_1_bits_26),
    .io_in_1_bits_27(dataIn_mux_io_in_1_bits_27),
    .io_in_1_bits_28(dataIn_mux_io_in_1_bits_28),
    .io_in_1_bits_29(dataIn_mux_io_in_1_bits_29),
    .io_in_1_bits_30(dataIn_mux_io_in_1_bits_30),
    .io_in_1_bits_31(dataIn_mux_io_in_1_bits_31),
    .io_sel_ready(dataIn_mux_io_sel_ready),
    .io_sel_valid(dataIn_mux_io_sel_valid),
    .io_sel_bits(dataIn_mux_io_sel_bits),
    .io_out_ready(dataIn_mux_io_out_ready),
    .io_out_valid(dataIn_mux_io_out_valid),
    .io_out_bits_0(dataIn_mux_io_out_bits_0),
    .io_out_bits_1(dataIn_mux_io_out_bits_1),
    .io_out_bits_2(dataIn_mux_io_out_bits_2),
    .io_out_bits_3(dataIn_mux_io_out_bits_3),
    .io_out_bits_4(dataIn_mux_io_out_bits_4),
    .io_out_bits_5(dataIn_mux_io_out_bits_5),
    .io_out_bits_6(dataIn_mux_io_out_bits_6),
    .io_out_bits_7(dataIn_mux_io_out_bits_7),
    .io_out_bits_8(dataIn_mux_io_out_bits_8),
    .io_out_bits_9(dataIn_mux_io_out_bits_9),
    .io_out_bits_10(dataIn_mux_io_out_bits_10),
    .io_out_bits_11(dataIn_mux_io_out_bits_11),
    .io_out_bits_12(dataIn_mux_io_out_bits_12),
    .io_out_bits_13(dataIn_mux_io_out_bits_13),
    .io_out_bits_14(dataIn_mux_io_out_bits_14),
    .io_out_bits_15(dataIn_mux_io_out_bits_15),
    .io_out_bits_16(dataIn_mux_io_out_bits_16),
    .io_out_bits_17(dataIn_mux_io_out_bits_17),
    .io_out_bits_18(dataIn_mux_io_out_bits_18),
    .io_out_bits_19(dataIn_mux_io_out_bits_19),
    .io_out_bits_20(dataIn_mux_io_out_bits_20),
    .io_out_bits_21(dataIn_mux_io_out_bits_21),
    .io_out_bits_22(dataIn_mux_io_out_bits_22),
    .io_out_bits_23(dataIn_mux_io_out_bits_23),
    .io_out_bits_24(dataIn_mux_io_out_bits_24),
    .io_out_bits_25(dataIn_mux_io_out_bits_25),
    .io_out_bits_26(dataIn_mux_io_out_bits_26),
    .io_out_bits_27(dataIn_mux_io_out_bits_27),
    .io_out_bits_28(dataIn_mux_io_out_bits_28),
    .io_out_bits_29(dataIn_mux_io_out_bits_29),
    .io_out_bits_30(dataIn_mux_io_out_bits_30),
    .io_out_bits_31(dataIn_mux_io_out_bits_31)
  );
  Demux dataOut_demux ( // @[Demux.scala 46:23]
    .io_in_ready(dataOut_demux_io_in_ready),
    .io_in_valid(dataOut_demux_io_in_valid),
    .io_in_bits_0(dataOut_demux_io_in_bits_0),
    .io_in_bits_1(dataOut_demux_io_in_bits_1),
    .io_in_bits_2(dataOut_demux_io_in_bits_2),
    .io_in_bits_3(dataOut_demux_io_in_bits_3),
    .io_in_bits_4(dataOut_demux_io_in_bits_4),
    .io_in_bits_5(dataOut_demux_io_in_bits_5),
    .io_in_bits_6(dataOut_demux_io_in_bits_6),
    .io_in_bits_7(dataOut_demux_io_in_bits_7),
    .io_in_bits_8(dataOut_demux_io_in_bits_8),
    .io_in_bits_9(dataOut_demux_io_in_bits_9),
    .io_in_bits_10(dataOut_demux_io_in_bits_10),
    .io_in_bits_11(dataOut_demux_io_in_bits_11),
    .io_in_bits_12(dataOut_demux_io_in_bits_12),
    .io_in_bits_13(dataOut_demux_io_in_bits_13),
    .io_in_bits_14(dataOut_demux_io_in_bits_14),
    .io_in_bits_15(dataOut_demux_io_in_bits_15),
    .io_in_bits_16(dataOut_demux_io_in_bits_16),
    .io_in_bits_17(dataOut_demux_io_in_bits_17),
    .io_in_bits_18(dataOut_demux_io_in_bits_18),
    .io_in_bits_19(dataOut_demux_io_in_bits_19),
    .io_in_bits_20(dataOut_demux_io_in_bits_20),
    .io_in_bits_21(dataOut_demux_io_in_bits_21),
    .io_in_bits_22(dataOut_demux_io_in_bits_22),
    .io_in_bits_23(dataOut_demux_io_in_bits_23),
    .io_in_bits_24(dataOut_demux_io_in_bits_24),
    .io_in_bits_25(dataOut_demux_io_in_bits_25),
    .io_in_bits_26(dataOut_demux_io_in_bits_26),
    .io_in_bits_27(dataOut_demux_io_in_bits_27),
    .io_in_bits_28(dataOut_demux_io_in_bits_28),
    .io_in_bits_29(dataOut_demux_io_in_bits_29),
    .io_in_bits_30(dataOut_demux_io_in_bits_30),
    .io_in_bits_31(dataOut_demux_io_in_bits_31),
    .io_sel_ready(dataOut_demux_io_sel_ready),
    .io_sel_valid(dataOut_demux_io_sel_valid),
    .io_sel_bits(dataOut_demux_io_sel_bits),
    .io_out_0_ready(dataOut_demux_io_out_0_ready),
    .io_out_0_valid(dataOut_demux_io_out_0_valid),
    .io_out_0_bits_0(dataOut_demux_io_out_0_bits_0),
    .io_out_0_bits_1(dataOut_demux_io_out_0_bits_1),
    .io_out_0_bits_2(dataOut_demux_io_out_0_bits_2),
    .io_out_0_bits_3(dataOut_demux_io_out_0_bits_3),
    .io_out_0_bits_4(dataOut_demux_io_out_0_bits_4),
    .io_out_0_bits_5(dataOut_demux_io_out_0_bits_5),
    .io_out_0_bits_6(dataOut_demux_io_out_0_bits_6),
    .io_out_0_bits_7(dataOut_demux_io_out_0_bits_7),
    .io_out_0_bits_8(dataOut_demux_io_out_0_bits_8),
    .io_out_0_bits_9(dataOut_demux_io_out_0_bits_9),
    .io_out_0_bits_10(dataOut_demux_io_out_0_bits_10),
    .io_out_0_bits_11(dataOut_demux_io_out_0_bits_11),
    .io_out_0_bits_12(dataOut_demux_io_out_0_bits_12),
    .io_out_0_bits_13(dataOut_demux_io_out_0_bits_13),
    .io_out_0_bits_14(dataOut_demux_io_out_0_bits_14),
    .io_out_0_bits_15(dataOut_demux_io_out_0_bits_15),
    .io_out_0_bits_16(dataOut_demux_io_out_0_bits_16),
    .io_out_0_bits_17(dataOut_demux_io_out_0_bits_17),
    .io_out_0_bits_18(dataOut_demux_io_out_0_bits_18),
    .io_out_0_bits_19(dataOut_demux_io_out_0_bits_19),
    .io_out_0_bits_20(dataOut_demux_io_out_0_bits_20),
    .io_out_0_bits_21(dataOut_demux_io_out_0_bits_21),
    .io_out_0_bits_22(dataOut_demux_io_out_0_bits_22),
    .io_out_0_bits_23(dataOut_demux_io_out_0_bits_23),
    .io_out_0_bits_24(dataOut_demux_io_out_0_bits_24),
    .io_out_0_bits_25(dataOut_demux_io_out_0_bits_25),
    .io_out_0_bits_26(dataOut_demux_io_out_0_bits_26),
    .io_out_0_bits_27(dataOut_demux_io_out_0_bits_27),
    .io_out_0_bits_28(dataOut_demux_io_out_0_bits_28),
    .io_out_0_bits_29(dataOut_demux_io_out_0_bits_29),
    .io_out_0_bits_30(dataOut_demux_io_out_0_bits_30),
    .io_out_0_bits_31(dataOut_demux_io_out_0_bits_31),
    .io_out_1_ready(dataOut_demux_io_out_1_ready),
    .io_out_1_valid(dataOut_demux_io_out_1_valid),
    .io_out_1_bits_0(dataOut_demux_io_out_1_bits_0),
    .io_out_1_bits_1(dataOut_demux_io_out_1_bits_1),
    .io_out_1_bits_2(dataOut_demux_io_out_1_bits_2),
    .io_out_1_bits_3(dataOut_demux_io_out_1_bits_3),
    .io_out_1_bits_4(dataOut_demux_io_out_1_bits_4),
    .io_out_1_bits_5(dataOut_demux_io_out_1_bits_5),
    .io_out_1_bits_6(dataOut_demux_io_out_1_bits_6),
    .io_out_1_bits_7(dataOut_demux_io_out_1_bits_7),
    .io_out_1_bits_8(dataOut_demux_io_out_1_bits_8),
    .io_out_1_bits_9(dataOut_demux_io_out_1_bits_9),
    .io_out_1_bits_10(dataOut_demux_io_out_1_bits_10),
    .io_out_1_bits_11(dataOut_demux_io_out_1_bits_11),
    .io_out_1_bits_12(dataOut_demux_io_out_1_bits_12),
    .io_out_1_bits_13(dataOut_demux_io_out_1_bits_13),
    .io_out_1_bits_14(dataOut_demux_io_out_1_bits_14),
    .io_out_1_bits_15(dataOut_demux_io_out_1_bits_15),
    .io_out_1_bits_16(dataOut_demux_io_out_1_bits_16),
    .io_out_1_bits_17(dataOut_demux_io_out_1_bits_17),
    .io_out_1_bits_18(dataOut_demux_io_out_1_bits_18),
    .io_out_1_bits_19(dataOut_demux_io_out_1_bits_19),
    .io_out_1_bits_20(dataOut_demux_io_out_1_bits_20),
    .io_out_1_bits_21(dataOut_demux_io_out_1_bits_21),
    .io_out_1_bits_22(dataOut_demux_io_out_1_bits_22),
    .io_out_1_bits_23(dataOut_demux_io_out_1_bits_23),
    .io_out_1_bits_24(dataOut_demux_io_out_1_bits_24),
    .io_out_1_bits_25(dataOut_demux_io_out_1_bits_25),
    .io_out_1_bits_26(dataOut_demux_io_out_1_bits_26),
    .io_out_1_bits_27(dataOut_demux_io_out_1_bits_27),
    .io_out_1_bits_28(dataOut_demux_io_out_1_bits_28),
    .io_out_1_bits_29(dataOut_demux_io_out_1_bits_29),
    .io_out_1_bits_30(dataOut_demux_io_out_1_bits_30),
    .io_out_1_bits_31(dataOut_demux_io_out_1_bits_31)
  );
  assign io_control_ready = isDataIn & dataIn_mux_io_sel_ready | isDataOut & dataOut_demux_io_sel_ready; // @[HostRouter.scala 41:47]
  assign io_dram0_dataIn_ready = dataIn_mux_io_in_0_ready; // @[Mux.scala 79:18]
  assign io_dram0_dataOut_valid = dataOut_demux_io_out_0_valid; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_0 = dataOut_demux_io_out_0_bits_0; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_1 = dataOut_demux_io_out_0_bits_1; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_2 = dataOut_demux_io_out_0_bits_2; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_3 = dataOut_demux_io_out_0_bits_3; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_4 = dataOut_demux_io_out_0_bits_4; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_5 = dataOut_demux_io_out_0_bits_5; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_6 = dataOut_demux_io_out_0_bits_6; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_7 = dataOut_demux_io_out_0_bits_7; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_8 = dataOut_demux_io_out_0_bits_8; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_9 = dataOut_demux_io_out_0_bits_9; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_10 = dataOut_demux_io_out_0_bits_10; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_11 = dataOut_demux_io_out_0_bits_11; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_12 = dataOut_demux_io_out_0_bits_12; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_13 = dataOut_demux_io_out_0_bits_13; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_14 = dataOut_demux_io_out_0_bits_14; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_15 = dataOut_demux_io_out_0_bits_15; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_16 = dataOut_demux_io_out_0_bits_16; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_17 = dataOut_demux_io_out_0_bits_17; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_18 = dataOut_demux_io_out_0_bits_18; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_19 = dataOut_demux_io_out_0_bits_19; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_20 = dataOut_demux_io_out_0_bits_20; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_21 = dataOut_demux_io_out_0_bits_21; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_22 = dataOut_demux_io_out_0_bits_22; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_23 = dataOut_demux_io_out_0_bits_23; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_24 = dataOut_demux_io_out_0_bits_24; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_25 = dataOut_demux_io_out_0_bits_25; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_26 = dataOut_demux_io_out_0_bits_26; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_27 = dataOut_demux_io_out_0_bits_27; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_28 = dataOut_demux_io_out_0_bits_28; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_29 = dataOut_demux_io_out_0_bits_29; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_30 = dataOut_demux_io_out_0_bits_30; // @[Demux.scala 55:10]
  assign io_dram0_dataOut_bits_31 = dataOut_demux_io_out_0_bits_31; // @[Demux.scala 55:10]
  assign io_dram1_dataIn_ready = dataIn_mux_io_in_1_ready; // @[Mux.scala 80:18]
  assign io_dram1_dataOut_valid = dataOut_demux_io_out_1_valid; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_0 = dataOut_demux_io_out_1_bits_0; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_1 = dataOut_demux_io_out_1_bits_1; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_2 = dataOut_demux_io_out_1_bits_2; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_3 = dataOut_demux_io_out_1_bits_3; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_4 = dataOut_demux_io_out_1_bits_4; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_5 = dataOut_demux_io_out_1_bits_5; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_6 = dataOut_demux_io_out_1_bits_6; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_7 = dataOut_demux_io_out_1_bits_7; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_8 = dataOut_demux_io_out_1_bits_8; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_9 = dataOut_demux_io_out_1_bits_9; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_10 = dataOut_demux_io_out_1_bits_10; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_11 = dataOut_demux_io_out_1_bits_11; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_12 = dataOut_demux_io_out_1_bits_12; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_13 = dataOut_demux_io_out_1_bits_13; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_14 = dataOut_demux_io_out_1_bits_14; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_15 = dataOut_demux_io_out_1_bits_15; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_16 = dataOut_demux_io_out_1_bits_16; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_17 = dataOut_demux_io_out_1_bits_17; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_18 = dataOut_demux_io_out_1_bits_18; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_19 = dataOut_demux_io_out_1_bits_19; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_20 = dataOut_demux_io_out_1_bits_20; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_21 = dataOut_demux_io_out_1_bits_21; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_22 = dataOut_demux_io_out_1_bits_22; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_23 = dataOut_demux_io_out_1_bits_23; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_24 = dataOut_demux_io_out_1_bits_24; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_25 = dataOut_demux_io_out_1_bits_25; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_26 = dataOut_demux_io_out_1_bits_26; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_27 = dataOut_demux_io_out_1_bits_27; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_28 = dataOut_demux_io_out_1_bits_28; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_29 = dataOut_demux_io_out_1_bits_29; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_30 = dataOut_demux_io_out_1_bits_30; // @[Demux.scala 56:10]
  assign io_dram1_dataOut_bits_31 = dataOut_demux_io_out_1_bits_31; // @[Demux.scala 56:10]
  assign io_mem_output_ready = dataOut_demux_io_in_ready; // @[Demux.scala 54:17]
  assign io_mem_input_valid = dataIn_mux_io_out_valid; // @[Mux.scala 81:9]
  assign io_mem_input_bits_0 = dataIn_mux_io_out_bits_0; // @[Mux.scala 81:9]
  assign io_mem_input_bits_1 = dataIn_mux_io_out_bits_1; // @[Mux.scala 81:9]
  assign io_mem_input_bits_2 = dataIn_mux_io_out_bits_2; // @[Mux.scala 81:9]
  assign io_mem_input_bits_3 = dataIn_mux_io_out_bits_3; // @[Mux.scala 81:9]
  assign io_mem_input_bits_4 = dataIn_mux_io_out_bits_4; // @[Mux.scala 81:9]
  assign io_mem_input_bits_5 = dataIn_mux_io_out_bits_5; // @[Mux.scala 81:9]
  assign io_mem_input_bits_6 = dataIn_mux_io_out_bits_6; // @[Mux.scala 81:9]
  assign io_mem_input_bits_7 = dataIn_mux_io_out_bits_7; // @[Mux.scala 81:9]
  assign io_mem_input_bits_8 = dataIn_mux_io_out_bits_8; // @[Mux.scala 81:9]
  assign io_mem_input_bits_9 = dataIn_mux_io_out_bits_9; // @[Mux.scala 81:9]
  assign io_mem_input_bits_10 = dataIn_mux_io_out_bits_10; // @[Mux.scala 81:9]
  assign io_mem_input_bits_11 = dataIn_mux_io_out_bits_11; // @[Mux.scala 81:9]
  assign io_mem_input_bits_12 = dataIn_mux_io_out_bits_12; // @[Mux.scala 81:9]
  assign io_mem_input_bits_13 = dataIn_mux_io_out_bits_13; // @[Mux.scala 81:9]
  assign io_mem_input_bits_14 = dataIn_mux_io_out_bits_14; // @[Mux.scala 81:9]
  assign io_mem_input_bits_15 = dataIn_mux_io_out_bits_15; // @[Mux.scala 81:9]
  assign io_mem_input_bits_16 = dataIn_mux_io_out_bits_16; // @[Mux.scala 81:9]
  assign io_mem_input_bits_17 = dataIn_mux_io_out_bits_17; // @[Mux.scala 81:9]
  assign io_mem_input_bits_18 = dataIn_mux_io_out_bits_18; // @[Mux.scala 81:9]
  assign io_mem_input_bits_19 = dataIn_mux_io_out_bits_19; // @[Mux.scala 81:9]
  assign io_mem_input_bits_20 = dataIn_mux_io_out_bits_20; // @[Mux.scala 81:9]
  assign io_mem_input_bits_21 = dataIn_mux_io_out_bits_21; // @[Mux.scala 81:9]
  assign io_mem_input_bits_22 = dataIn_mux_io_out_bits_22; // @[Mux.scala 81:9]
  assign io_mem_input_bits_23 = dataIn_mux_io_out_bits_23; // @[Mux.scala 81:9]
  assign io_mem_input_bits_24 = dataIn_mux_io_out_bits_24; // @[Mux.scala 81:9]
  assign io_mem_input_bits_25 = dataIn_mux_io_out_bits_25; // @[Mux.scala 81:9]
  assign io_mem_input_bits_26 = dataIn_mux_io_out_bits_26; // @[Mux.scala 81:9]
  assign io_mem_input_bits_27 = dataIn_mux_io_out_bits_27; // @[Mux.scala 81:9]
  assign io_mem_input_bits_28 = dataIn_mux_io_out_bits_28; // @[Mux.scala 81:9]
  assign io_mem_input_bits_29 = dataIn_mux_io_out_bits_29; // @[Mux.scala 81:9]
  assign io_mem_input_bits_30 = dataIn_mux_io_out_bits_30; // @[Mux.scala 81:9]
  assign io_mem_input_bits_31 = dataIn_mux_io_out_bits_31; // @[Mux.scala 81:9]
  assign dataIn_mux_io_in_0_valid = io_dram0_dataIn_valid; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_0 = io_dram0_dataIn_bits_0; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_1 = io_dram0_dataIn_bits_1; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_2 = io_dram0_dataIn_bits_2; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_3 = io_dram0_dataIn_bits_3; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_4 = io_dram0_dataIn_bits_4; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_5 = io_dram0_dataIn_bits_5; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_6 = io_dram0_dataIn_bits_6; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_7 = io_dram0_dataIn_bits_7; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_8 = io_dram0_dataIn_bits_8; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_9 = io_dram0_dataIn_bits_9; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_10 = io_dram0_dataIn_bits_10; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_11 = io_dram0_dataIn_bits_11; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_12 = io_dram0_dataIn_bits_12; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_13 = io_dram0_dataIn_bits_13; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_14 = io_dram0_dataIn_bits_14; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_15 = io_dram0_dataIn_bits_15; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_16 = io_dram0_dataIn_bits_16; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_17 = io_dram0_dataIn_bits_17; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_18 = io_dram0_dataIn_bits_18; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_19 = io_dram0_dataIn_bits_19; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_20 = io_dram0_dataIn_bits_20; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_21 = io_dram0_dataIn_bits_21; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_22 = io_dram0_dataIn_bits_22; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_23 = io_dram0_dataIn_bits_23; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_24 = io_dram0_dataIn_bits_24; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_25 = io_dram0_dataIn_bits_25; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_26 = io_dram0_dataIn_bits_26; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_27 = io_dram0_dataIn_bits_27; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_28 = io_dram0_dataIn_bits_28; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_29 = io_dram0_dataIn_bits_29; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_30 = io_dram0_dataIn_bits_30; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_0_bits_31 = io_dram0_dataIn_bits_31; // @[Mux.scala 79:18]
  assign dataIn_mux_io_in_1_valid = io_dram1_dataIn_valid; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_0 = io_dram1_dataIn_bits_0; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_1 = io_dram1_dataIn_bits_1; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_2 = io_dram1_dataIn_bits_2; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_3 = io_dram1_dataIn_bits_3; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_4 = io_dram1_dataIn_bits_4; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_5 = io_dram1_dataIn_bits_5; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_6 = io_dram1_dataIn_bits_6; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_7 = io_dram1_dataIn_bits_7; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_8 = io_dram1_dataIn_bits_8; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_9 = io_dram1_dataIn_bits_9; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_10 = io_dram1_dataIn_bits_10; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_11 = io_dram1_dataIn_bits_11; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_12 = io_dram1_dataIn_bits_12; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_13 = io_dram1_dataIn_bits_13; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_14 = io_dram1_dataIn_bits_14; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_15 = io_dram1_dataIn_bits_15; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_16 = io_dram1_dataIn_bits_16; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_17 = io_dram1_dataIn_bits_17; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_18 = io_dram1_dataIn_bits_18; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_19 = io_dram1_dataIn_bits_19; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_20 = io_dram1_dataIn_bits_20; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_21 = io_dram1_dataIn_bits_21; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_22 = io_dram1_dataIn_bits_22; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_23 = io_dram1_dataIn_bits_23; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_24 = io_dram1_dataIn_bits_24; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_25 = io_dram1_dataIn_bits_25; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_26 = io_dram1_dataIn_bits_26; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_27 = io_dram1_dataIn_bits_27; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_28 = io_dram1_dataIn_bits_28; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_29 = io_dram1_dataIn_bits_29; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_30 = io_dram1_dataIn_bits_30; // @[Mux.scala 80:18]
  assign dataIn_mux_io_in_1_bits_31 = io_dram1_dataIn_bits_31; // @[Mux.scala 80:18]
  assign dataIn_mux_io_sel_valid = io_control_valid & isDataIn; // @[HostRouter.scala 43:33]
  assign dataIn_mux_io_sel_bits = io_control_bits_kind[1]; // @[HostRouter.scala 44:35]
  assign dataIn_mux_io_out_ready = io_mem_input_ready; // @[Mux.scala 81:9]
  assign dataOut_demux_io_in_valid = io_mem_output_valid; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_0 = io_mem_output_bits_0; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_1 = io_mem_output_bits_1; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_2 = io_mem_output_bits_2; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_3 = io_mem_output_bits_3; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_4 = io_mem_output_bits_4; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_5 = io_mem_output_bits_5; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_6 = io_mem_output_bits_6; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_7 = io_mem_output_bits_7; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_8 = io_mem_output_bits_8; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_9 = io_mem_output_bits_9; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_10 = io_mem_output_bits_10; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_11 = io_mem_output_bits_11; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_12 = io_mem_output_bits_12; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_13 = io_mem_output_bits_13; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_14 = io_mem_output_bits_14; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_15 = io_mem_output_bits_15; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_16 = io_mem_output_bits_16; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_17 = io_mem_output_bits_17; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_18 = io_mem_output_bits_18; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_19 = io_mem_output_bits_19; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_20 = io_mem_output_bits_20; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_21 = io_mem_output_bits_21; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_22 = io_mem_output_bits_22; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_23 = io_mem_output_bits_23; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_24 = io_mem_output_bits_24; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_25 = io_mem_output_bits_25; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_26 = io_mem_output_bits_26; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_27 = io_mem_output_bits_27; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_28 = io_mem_output_bits_28; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_29 = io_mem_output_bits_29; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_30 = io_mem_output_bits_30; // @[Demux.scala 54:17]
  assign dataOut_demux_io_in_bits_31 = io_mem_output_bits_31; // @[Demux.scala 54:17]
  assign dataOut_demux_io_sel_valid = io_control_valid & isDataOut; // @[HostRouter.scala 46:34]
  assign dataOut_demux_io_sel_bits = io_control_bits_kind[1]; // @[HostRouter.scala 47:36]
  assign dataOut_demux_io_out_0_ready = io_dram0_dataOut_ready; // @[Demux.scala 55:10]
  assign dataOut_demux_io_out_1_ready = io_dram1_dataOut_ready; // @[Demux.scala 56:10]
endmodule
module Queue_28(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_instruction_op,
  input         io_enq_bits_instruction_sourceLeft,
  input         io_enq_bits_instruction_sourceRight,
  input         io_enq_bits_instruction_dest,
  input  [11:0] io_enq_bits_readAddress,
  input  [11:0] io_enq_bits_writeAddress,
  input         io_enq_bits_accumulate,
  input         io_enq_bits_write,
  input         io_enq_bits_read,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_instruction_op,
  output        io_deq_bits_instruction_sourceLeft,
  output        io_deq_bits_instruction_sourceRight,
  output        io_deq_bits_instruction_dest,
  output [11:0] io_deq_bits_readAddress,
  output [11:0] io_deq_bits_writeAddress,
  output        io_deq_bits_accumulate,
  output        io_deq_bits_write,
  output        io_deq_bits_read
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_instruction_op [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_instruction_op_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_instruction_op_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_instruction_op_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_instruction_op_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_instruction_op_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_op_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_instruction_op_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_instruction_sourceLeft [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceLeft_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_instruction_sourceRight [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_instruction_sourceRight_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_instruction_dest [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_instruction_dest_MPORT_en; // @[Decoupled.scala 259:95]
  reg [11:0] ram_readAddress [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_readAddress_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_readAddress_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [11:0] ram_readAddress_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [11:0] ram_readAddress_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_readAddress_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_readAddress_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_readAddress_MPORT_en; // @[Decoupled.scala 259:95]
  reg [11:0] ram_writeAddress [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_writeAddress_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_writeAddress_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [11:0] ram_writeAddress_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [11:0] ram_writeAddress_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_writeAddress_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_writeAddress_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_writeAddress_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_accumulate [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_accumulate_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_write [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_read [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_read_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_read_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_read_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_en; // @[Decoupled.scala 259:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_instruction_op_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instruction_op_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instruction_op_io_deq_bits_MPORT_data = ram_instruction_op[ram_instruction_op_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_instruction_op_MPORT_data = io_enq_bits_instruction_op;
  assign ram_instruction_op_MPORT_addr = enq_ptr_value;
  assign ram_instruction_op_MPORT_mask = 1'h1;
  assign ram_instruction_op_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_instruction_sourceLeft_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instruction_sourceLeft_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instruction_sourceLeft_io_deq_bits_MPORT_data =
    ram_instruction_sourceLeft[ram_instruction_sourceLeft_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_instruction_sourceLeft_MPORT_data = io_enq_bits_instruction_sourceLeft;
  assign ram_instruction_sourceLeft_MPORT_addr = enq_ptr_value;
  assign ram_instruction_sourceLeft_MPORT_mask = 1'h1;
  assign ram_instruction_sourceLeft_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_instruction_sourceRight_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instruction_sourceRight_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instruction_sourceRight_io_deq_bits_MPORT_data =
    ram_instruction_sourceRight[ram_instruction_sourceRight_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_instruction_sourceRight_MPORT_data = io_enq_bits_instruction_sourceRight;
  assign ram_instruction_sourceRight_MPORT_addr = enq_ptr_value;
  assign ram_instruction_sourceRight_MPORT_mask = 1'h1;
  assign ram_instruction_sourceRight_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_instruction_dest_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instruction_dest_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instruction_dest_io_deq_bits_MPORT_data = ram_instruction_dest[ram_instruction_dest_io_deq_bits_MPORT_addr]
    ; // @[Decoupled.scala 259:95]
  assign ram_instruction_dest_MPORT_data = io_enq_bits_instruction_dest;
  assign ram_instruction_dest_MPORT_addr = enq_ptr_value;
  assign ram_instruction_dest_MPORT_mask = 1'h1;
  assign ram_instruction_dest_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_readAddress_io_deq_bits_MPORT_en = 1'h1;
  assign ram_readAddress_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_readAddress_io_deq_bits_MPORT_data = ram_readAddress[ram_readAddress_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_readAddress_MPORT_data = io_enq_bits_readAddress;
  assign ram_readAddress_MPORT_addr = enq_ptr_value;
  assign ram_readAddress_MPORT_mask = 1'h1;
  assign ram_readAddress_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_writeAddress_io_deq_bits_MPORT_en = 1'h1;
  assign ram_writeAddress_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_writeAddress_io_deq_bits_MPORT_data = ram_writeAddress[ram_writeAddress_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_writeAddress_MPORT_data = io_enq_bits_writeAddress;
  assign ram_writeAddress_MPORT_addr = enq_ptr_value;
  assign ram_writeAddress_MPORT_mask = 1'h1;
  assign ram_writeAddress_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_accumulate_io_deq_bits_MPORT_en = 1'h1;
  assign ram_accumulate_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_accumulate_io_deq_bits_MPORT_data = ram_accumulate[ram_accumulate_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_accumulate_MPORT_data = io_enq_bits_accumulate;
  assign ram_accumulate_MPORT_addr = enq_ptr_value;
  assign ram_accumulate_MPORT_mask = 1'h1;
  assign ram_accumulate_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_write_io_deq_bits_MPORT_en = 1'h1;
  assign ram_write_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_write_io_deq_bits_MPORT_data = ram_write[ram_write_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_write_MPORT_data = io_enq_bits_write;
  assign ram_write_MPORT_addr = enq_ptr_value;
  assign ram_write_MPORT_mask = 1'h1;
  assign ram_write_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_read_io_deq_bits_MPORT_en = 1'h1;
  assign ram_read_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_read_io_deq_bits_MPORT_data = ram_read[ram_read_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_read_MPORT_data = io_enq_bits_read;
  assign ram_read_MPORT_addr = enq_ptr_value;
  assign ram_read_MPORT_mask = 1'h1;
  assign ram_read_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_instruction_op = ram_instruction_op_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_instruction_sourceLeft = ram_instruction_sourceLeft_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_instruction_sourceRight = ram_instruction_sourceRight_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_instruction_dest = ram_instruction_dest_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_readAddress = ram_readAddress_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_writeAddress = ram_writeAddress_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_accumulate = ram_accumulate_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_write = ram_write_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_read = ram_read_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_instruction_op_MPORT_en & ram_instruction_op_MPORT_mask) begin
      ram_instruction_op[ram_instruction_op_MPORT_addr] <= ram_instruction_op_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_instruction_sourceLeft_MPORT_en & ram_instruction_sourceLeft_MPORT_mask) begin
      ram_instruction_sourceLeft[ram_instruction_sourceLeft_MPORT_addr] <= ram_instruction_sourceLeft_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_instruction_sourceRight_MPORT_en & ram_instruction_sourceRight_MPORT_mask) begin
      ram_instruction_sourceRight[ram_instruction_sourceRight_MPORT_addr] <= ram_instruction_sourceRight_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_instruction_dest_MPORT_en & ram_instruction_dest_MPORT_mask) begin
      ram_instruction_dest[ram_instruction_dest_MPORT_addr] <= ram_instruction_dest_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_readAddress_MPORT_en & ram_readAddress_MPORT_mask) begin
      ram_readAddress[ram_readAddress_MPORT_addr] <= ram_readAddress_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_writeAddress_MPORT_en & ram_writeAddress_MPORT_mask) begin
      ram_writeAddress[ram_writeAddress_MPORT_addr] <= ram_writeAddress_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_accumulate_MPORT_en & ram_accumulate_MPORT_mask) begin
      ram_accumulate[ram_accumulate_MPORT_addr] <= ram_accumulate_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_write_MPORT_en & ram_write_MPORT_mask) begin
      ram_write[ram_write_MPORT_addr] <= ram_write_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_read_MPORT_en & ram_read_MPORT_mask) begin
      ram_read[ram_read_MPORT_addr] <= ram_read_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_instruction_op[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_instruction_sourceLeft[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_instruction_sourceRight[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_instruction_dest[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_readAddress[initvar] = _RAND_4[11:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_writeAddress[initvar] = _RAND_5[11:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_accumulate[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_write[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_read[initvar] = _RAND_8[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  enq_ptr_value = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  deq_ptr_value = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  maybe_full = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_29(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_load,
  input   io_enq_bits_zeroes,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits_load,
  output  io_deq_bits_zeroes
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  ram_load [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_load_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_load_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_load_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_load_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_load_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_load_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_load_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_zeroes [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_zeroes_MPORT_en; // @[Decoupled.scala 259:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_load_io_deq_bits_MPORT_en = 1'h1;
  assign ram_load_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_load_io_deq_bits_MPORT_data = ram_load[ram_load_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_load_MPORT_data = io_enq_bits_load;
  assign ram_load_MPORT_addr = enq_ptr_value;
  assign ram_load_MPORT_mask = 1'h1;
  assign ram_load_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_zeroes_io_deq_bits_MPORT_en = 1'h1;
  assign ram_zeroes_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_zeroes_io_deq_bits_MPORT_data = ram_zeroes[ram_zeroes_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_zeroes_MPORT_data = io_enq_bits_zeroes;
  assign ram_zeroes_MPORT_addr = enq_ptr_value;
  assign ram_zeroes_MPORT_mask = 1'h1;
  assign ram_zeroes_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_load = ram_load_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_zeroes = ram_zeroes_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_load_MPORT_en & ram_load_MPORT_mask) begin
      ram_load[ram_load_MPORT_addr] <= ram_load_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_zeroes_MPORT_en & ram_zeroes_MPORT_mask) begin
      ram_zeroes[ram_zeroes_MPORT_addr] <= ram_zeroes_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_load[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_zeroes[initvar] = _RAND_1[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TCU(
  input         clock,
  input         reset,
  output        io_instruction_ready,
  input         io_instruction_valid,
  input  [3:0]  io_instruction_bits_opcode,
  input  [3:0]  io_instruction_bits_flags,
  input  [63:0] io_instruction_bits_arguments,
  input         io_dram0_control_ready,
  output        io_dram0_control_valid,
  output        io_dram0_control_bits_write,
  output [20:0] io_dram0_control_bits_address,
  output [20:0] io_dram0_control_bits_size,
  output        io_dram0_dataIn_ready,
  input         io_dram0_dataIn_valid,
  input  [15:0] io_dram0_dataIn_bits_0,
  input  [15:0] io_dram0_dataIn_bits_1,
  input  [15:0] io_dram0_dataIn_bits_2,
  input  [15:0] io_dram0_dataIn_bits_3,
  input  [15:0] io_dram0_dataIn_bits_4,
  input  [15:0] io_dram0_dataIn_bits_5,
  input  [15:0] io_dram0_dataIn_bits_6,
  input  [15:0] io_dram0_dataIn_bits_7,
  input  [15:0] io_dram0_dataIn_bits_8,
  input  [15:0] io_dram0_dataIn_bits_9,
  input  [15:0] io_dram0_dataIn_bits_10,
  input  [15:0] io_dram0_dataIn_bits_11,
  input  [15:0] io_dram0_dataIn_bits_12,
  input  [15:0] io_dram0_dataIn_bits_13,
  input  [15:0] io_dram0_dataIn_bits_14,
  input  [15:0] io_dram0_dataIn_bits_15,
  input  [15:0] io_dram0_dataIn_bits_16,
  input  [15:0] io_dram0_dataIn_bits_17,
  input  [15:0] io_dram0_dataIn_bits_18,
  input  [15:0] io_dram0_dataIn_bits_19,
  input  [15:0] io_dram0_dataIn_bits_20,
  input  [15:0] io_dram0_dataIn_bits_21,
  input  [15:0] io_dram0_dataIn_bits_22,
  input  [15:0] io_dram0_dataIn_bits_23,
  input  [15:0] io_dram0_dataIn_bits_24,
  input  [15:0] io_dram0_dataIn_bits_25,
  input  [15:0] io_dram0_dataIn_bits_26,
  input  [15:0] io_dram0_dataIn_bits_27,
  input  [15:0] io_dram0_dataIn_bits_28,
  input  [15:0] io_dram0_dataIn_bits_29,
  input  [15:0] io_dram0_dataIn_bits_30,
  input  [15:0] io_dram0_dataIn_bits_31,
  input         io_dram0_dataOut_ready,
  output        io_dram0_dataOut_valid,
  output [15:0] io_dram0_dataOut_bits_0,
  output [15:0] io_dram0_dataOut_bits_1,
  output [15:0] io_dram0_dataOut_bits_2,
  output [15:0] io_dram0_dataOut_bits_3,
  output [15:0] io_dram0_dataOut_bits_4,
  output [15:0] io_dram0_dataOut_bits_5,
  output [15:0] io_dram0_dataOut_bits_6,
  output [15:0] io_dram0_dataOut_bits_7,
  output [15:0] io_dram0_dataOut_bits_8,
  output [15:0] io_dram0_dataOut_bits_9,
  output [15:0] io_dram0_dataOut_bits_10,
  output [15:0] io_dram0_dataOut_bits_11,
  output [15:0] io_dram0_dataOut_bits_12,
  output [15:0] io_dram0_dataOut_bits_13,
  output [15:0] io_dram0_dataOut_bits_14,
  output [15:0] io_dram0_dataOut_bits_15,
  output [15:0] io_dram0_dataOut_bits_16,
  output [15:0] io_dram0_dataOut_bits_17,
  output [15:0] io_dram0_dataOut_bits_18,
  output [15:0] io_dram0_dataOut_bits_19,
  output [15:0] io_dram0_dataOut_bits_20,
  output [15:0] io_dram0_dataOut_bits_21,
  output [15:0] io_dram0_dataOut_bits_22,
  output [15:0] io_dram0_dataOut_bits_23,
  output [15:0] io_dram0_dataOut_bits_24,
  output [15:0] io_dram0_dataOut_bits_25,
  output [15:0] io_dram0_dataOut_bits_26,
  output [15:0] io_dram0_dataOut_bits_27,
  output [15:0] io_dram0_dataOut_bits_28,
  output [15:0] io_dram0_dataOut_bits_29,
  output [15:0] io_dram0_dataOut_bits_30,
  output [15:0] io_dram0_dataOut_bits_31,
  input         io_dram1_control_ready,
  output        io_dram1_control_valid,
  output        io_dram1_control_bits_write,
  output [20:0] io_dram1_control_bits_address,
  output [20:0] io_dram1_control_bits_size,
  output        io_dram1_dataIn_ready,
  input         io_dram1_dataIn_valid,
  input  [15:0] io_dram1_dataIn_bits_0,
  input  [15:0] io_dram1_dataIn_bits_1,
  input  [15:0] io_dram1_dataIn_bits_2,
  input  [15:0] io_dram1_dataIn_bits_3,
  input  [15:0] io_dram1_dataIn_bits_4,
  input  [15:0] io_dram1_dataIn_bits_5,
  input  [15:0] io_dram1_dataIn_bits_6,
  input  [15:0] io_dram1_dataIn_bits_7,
  input  [15:0] io_dram1_dataIn_bits_8,
  input  [15:0] io_dram1_dataIn_bits_9,
  input  [15:0] io_dram1_dataIn_bits_10,
  input  [15:0] io_dram1_dataIn_bits_11,
  input  [15:0] io_dram1_dataIn_bits_12,
  input  [15:0] io_dram1_dataIn_bits_13,
  input  [15:0] io_dram1_dataIn_bits_14,
  input  [15:0] io_dram1_dataIn_bits_15,
  input  [15:0] io_dram1_dataIn_bits_16,
  input  [15:0] io_dram1_dataIn_bits_17,
  input  [15:0] io_dram1_dataIn_bits_18,
  input  [15:0] io_dram1_dataIn_bits_19,
  input  [15:0] io_dram1_dataIn_bits_20,
  input  [15:0] io_dram1_dataIn_bits_21,
  input  [15:0] io_dram1_dataIn_bits_22,
  input  [15:0] io_dram1_dataIn_bits_23,
  input  [15:0] io_dram1_dataIn_bits_24,
  input  [15:0] io_dram1_dataIn_bits_25,
  input  [15:0] io_dram1_dataIn_bits_26,
  input  [15:0] io_dram1_dataIn_bits_27,
  input  [15:0] io_dram1_dataIn_bits_28,
  input  [15:0] io_dram1_dataIn_bits_29,
  input  [15:0] io_dram1_dataIn_bits_30,
  input  [15:0] io_dram1_dataIn_bits_31,
  input         io_dram1_dataOut_ready,
  output        io_dram1_dataOut_valid,
  output [15:0] io_dram1_dataOut_bits_0,
  output [15:0] io_dram1_dataOut_bits_1,
  output [15:0] io_dram1_dataOut_bits_2,
  output [15:0] io_dram1_dataOut_bits_3,
  output [15:0] io_dram1_dataOut_bits_4,
  output [15:0] io_dram1_dataOut_bits_5,
  output [15:0] io_dram1_dataOut_bits_6,
  output [15:0] io_dram1_dataOut_bits_7,
  output [15:0] io_dram1_dataOut_bits_8,
  output [15:0] io_dram1_dataOut_bits_9,
  output [15:0] io_dram1_dataOut_bits_10,
  output [15:0] io_dram1_dataOut_bits_11,
  output [15:0] io_dram1_dataOut_bits_12,
  output [15:0] io_dram1_dataOut_bits_13,
  output [15:0] io_dram1_dataOut_bits_14,
  output [15:0] io_dram1_dataOut_bits_15,
  output [15:0] io_dram1_dataOut_bits_16,
  output [15:0] io_dram1_dataOut_bits_17,
  output [15:0] io_dram1_dataOut_bits_18,
  output [15:0] io_dram1_dataOut_bits_19,
  output [15:0] io_dram1_dataOut_bits_20,
  output [15:0] io_dram1_dataOut_bits_21,
  output [15:0] io_dram1_dataOut_bits_22,
  output [15:0] io_dram1_dataOut_bits_23,
  output [15:0] io_dram1_dataOut_bits_24,
  output [15:0] io_dram1_dataOut_bits_25,
  output [15:0] io_dram1_dataOut_bits_26,
  output [15:0] io_dram1_dataOut_bits_27,
  output [15:0] io_dram1_dataOut_bits_28,
  output [15:0] io_dram1_dataOut_bits_29,
  output [15:0] io_dram1_dataOut_bits_30,
  output [15:0] io_dram1_dataOut_bits_31,
  output [31:0] io_config_dram0AddressOffset,
  output [3:0]  io_config_dram0CacheBehaviour,
  output [31:0] io_config_dram1AddressOffset,
  output [3:0]  io_config_dram1CacheBehaviour,
  output        io_timeout,
  output        io_tracepoint,
  output [31:0] io_programCounter
);
  wire  decoder_clock; // @[TCU.scala 64:23]
  wire  decoder_reset; // @[TCU.scala 64:23]
  wire  decoder_io_instruction_ready; // @[TCU.scala 64:23]
  wire  decoder_io_instruction_valid; // @[TCU.scala 64:23]
  wire [3:0] decoder_io_instruction_bits_opcode; // @[TCU.scala 64:23]
  wire [3:0] decoder_io_instruction_bits_flags; // @[TCU.scala 64:23]
  wire [63:0] decoder_io_instruction_bits_arguments; // @[TCU.scala 64:23]
  wire  decoder_io_memPortA_ready; // @[TCU.scala 64:23]
  wire  decoder_io_memPortA_valid; // @[TCU.scala 64:23]
  wire  decoder_io_memPortA_bits_write; // @[TCU.scala 64:23]
  wire [13:0] decoder_io_memPortA_bits_address; // @[TCU.scala 64:23]
  wire  decoder_io_memPortB_ready; // @[TCU.scala 64:23]
  wire  decoder_io_memPortB_valid; // @[TCU.scala 64:23]
  wire  decoder_io_memPortB_bits_write; // @[TCU.scala 64:23]
  wire [13:0] decoder_io_memPortB_bits_address; // @[TCU.scala 64:23]
  wire  decoder_io_dram0_ready; // @[TCU.scala 64:23]
  wire  decoder_io_dram0_valid; // @[TCU.scala 64:23]
  wire  decoder_io_dram0_bits_write; // @[TCU.scala 64:23]
  wire [20:0] decoder_io_dram0_bits_address; // @[TCU.scala 64:23]
  wire [20:0] decoder_io_dram0_bits_size; // @[TCU.scala 64:23]
  wire  decoder_io_dram1_ready; // @[TCU.scala 64:23]
  wire  decoder_io_dram1_valid; // @[TCU.scala 64:23]
  wire  decoder_io_dram1_bits_write; // @[TCU.scala 64:23]
  wire [20:0] decoder_io_dram1_bits_address; // @[TCU.scala 64:23]
  wire [20:0] decoder_io_dram1_bits_size; // @[TCU.scala 64:23]
  wire  decoder_io_dataflow_ready; // @[TCU.scala 64:23]
  wire  decoder_io_dataflow_valid; // @[TCU.scala 64:23]
  wire [3:0] decoder_io_dataflow_bits_kind; // @[TCU.scala 64:23]
  wire [13:0] decoder_io_dataflow_bits_size; // @[TCU.scala 64:23]
  wire  decoder_io_hostDataflow_ready; // @[TCU.scala 64:23]
  wire  decoder_io_hostDataflow_valid; // @[TCU.scala 64:23]
  wire [1:0] decoder_io_hostDataflow_bits_kind; // @[TCU.scala 64:23]
  wire  decoder_io_acc_ready; // @[TCU.scala 64:23]
  wire  decoder_io_acc_valid; // @[TCU.scala 64:23]
  wire [3:0] decoder_io_acc_bits_instruction_op; // @[TCU.scala 64:23]
  wire  decoder_io_acc_bits_instruction_sourceLeft; // @[TCU.scala 64:23]
  wire  decoder_io_acc_bits_instruction_sourceRight; // @[TCU.scala 64:23]
  wire  decoder_io_acc_bits_instruction_dest; // @[TCU.scala 64:23]
  wire [11:0] decoder_io_acc_bits_readAddress; // @[TCU.scala 64:23]
  wire [11:0] decoder_io_acc_bits_writeAddress; // @[TCU.scala 64:23]
  wire  decoder_io_acc_bits_accumulate; // @[TCU.scala 64:23]
  wire  decoder_io_acc_bits_write; // @[TCU.scala 64:23]
  wire  decoder_io_acc_bits_read; // @[TCU.scala 64:23]
  wire  decoder_io_array_ready; // @[TCU.scala 64:23]
  wire  decoder_io_array_valid; // @[TCU.scala 64:23]
  wire  decoder_io_array_bits_load; // @[TCU.scala 64:23]
  wire  decoder_io_array_bits_zeroes; // @[TCU.scala 64:23]
  wire [31:0] decoder_io_config_dram0AddressOffset; // @[TCU.scala 64:23]
  wire [3:0] decoder_io_config_dram0CacheBehaviour; // @[TCU.scala 64:23]
  wire [31:0] decoder_io_config_dram1AddressOffset; // @[TCU.scala 64:23]
  wire [3:0] decoder_io_config_dram1CacheBehaviour; // @[TCU.scala 64:23]
  wire  decoder_io_timeout; // @[TCU.scala 64:23]
  wire  decoder_io_error; // @[TCU.scala 64:23]
  wire  decoder_io_tracepoint; // @[TCU.scala 64:23]
  wire [31:0] decoder_io_programCounter; // @[TCU.scala 64:23]
  wire  array_clock; // @[TCU.scala 65:21]
  wire  array_reset; // @[TCU.scala 65:21]
  wire  array_io_control_ready; // @[TCU.scala 65:21]
  wire  array_io_control_valid; // @[TCU.scala 65:21]
  wire  array_io_control_bits_load; // @[TCU.scala 65:21]
  wire  array_io_control_bits_zeroes; // @[TCU.scala 65:21]
  wire  array_io_input_ready; // @[TCU.scala 65:21]
  wire  array_io_input_valid; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_0; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_1; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_2; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_3; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_4; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_5; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_6; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_7; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_8; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_9; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_10; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_11; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_12; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_13; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_14; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_15; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_16; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_17; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_18; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_19; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_20; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_21; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_22; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_23; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_24; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_25; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_26; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_27; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_28; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_29; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_30; // @[TCU.scala 65:21]
  wire [15:0] array_io_input_bits_31; // @[TCU.scala 65:21]
  wire  array_io_weight_ready; // @[TCU.scala 65:21]
  wire  array_io_weight_valid; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_0; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_1; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_2; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_3; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_4; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_5; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_6; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_7; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_8; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_9; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_10; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_11; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_12; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_13; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_14; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_15; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_16; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_17; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_18; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_19; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_20; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_21; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_22; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_23; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_24; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_25; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_26; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_27; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_28; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_29; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_30; // @[TCU.scala 65:21]
  wire [15:0] array_io_weight_bits_31; // @[TCU.scala 65:21]
  wire  array_io_output_ready; // @[TCU.scala 65:21]
  wire  array_io_output_valid; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_0; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_1; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_2; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_3; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_4; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_5; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_6; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_7; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_8; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_9; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_10; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_11; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_12; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_13; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_14; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_15; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_16; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_17; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_18; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_19; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_20; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_21; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_22; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_23; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_24; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_25; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_26; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_27; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_28; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_29; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_30; // @[TCU.scala 65:21]
  wire [15:0] array_io_output_bits_31; // @[TCU.scala 65:21]
  wire  acc_clock; // @[TCU.scala 68:19]
  wire  acc_reset; // @[TCU.scala 68:19]
  wire  acc_io_input_ready; // @[TCU.scala 68:19]
  wire  acc_io_input_valid; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_0; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_1; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_2; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_3; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_4; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_5; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_6; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_7; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_8; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_9; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_10; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_11; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_12; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_13; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_14; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_15; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_16; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_17; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_18; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_19; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_20; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_21; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_22; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_23; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_24; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_25; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_26; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_27; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_28; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_29; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_30; // @[TCU.scala 68:19]
  wire [15:0] acc_io_input_bits_31; // @[TCU.scala 68:19]
  wire  acc_io_output_ready; // @[TCU.scala 68:19]
  wire  acc_io_output_valid; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_0; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_1; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_2; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_3; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_4; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_5; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_6; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_7; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_8; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_9; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_10; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_11; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_12; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_13; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_14; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_15; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_16; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_17; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_18; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_19; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_20; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_21; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_22; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_23; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_24; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_25; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_26; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_27; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_28; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_29; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_30; // @[TCU.scala 68:19]
  wire [15:0] acc_io_output_bits_31; // @[TCU.scala 68:19]
  wire  acc_io_control_ready; // @[TCU.scala 68:19]
  wire  acc_io_control_valid; // @[TCU.scala 68:19]
  wire [3:0] acc_io_control_bits_instruction_op; // @[TCU.scala 68:19]
  wire  acc_io_control_bits_instruction_sourceLeft; // @[TCU.scala 68:19]
  wire  acc_io_control_bits_instruction_sourceRight; // @[TCU.scala 68:19]
  wire  acc_io_control_bits_instruction_dest; // @[TCU.scala 68:19]
  wire [11:0] acc_io_control_bits_readAddress; // @[TCU.scala 68:19]
  wire [11:0] acc_io_control_bits_writeAddress; // @[TCU.scala 68:19]
  wire  acc_io_control_bits_accumulate; // @[TCU.scala 68:19]
  wire  acc_io_control_bits_write; // @[TCU.scala 68:19]
  wire  acc_io_control_bits_read; // @[TCU.scala 68:19]
  wire  acc_io_tracepoint; // @[TCU.scala 68:19]
  wire [31:0] acc_io_programCounter; // @[TCU.scala 68:19]
  wire  mem_clock; // @[TCU.scala 71:19]
  wire  mem_reset; // @[TCU.scala 71:19]
  wire  mem_io_portA_control_ready; // @[TCU.scala 71:19]
  wire  mem_io_portA_control_valid; // @[TCU.scala 71:19]
  wire  mem_io_portA_control_bits_write; // @[TCU.scala 71:19]
  wire [13:0] mem_io_portA_control_bits_address; // @[TCU.scala 71:19]
  wire  mem_io_portA_input_ready; // @[TCU.scala 71:19]
  wire  mem_io_portA_input_valid; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_0; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_1; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_2; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_3; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_4; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_5; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_6; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_7; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_8; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_9; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_10; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_11; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_12; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_13; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_14; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_15; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_16; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_17; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_18; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_19; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_20; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_21; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_22; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_23; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_24; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_25; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_26; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_27; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_28; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_29; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_30; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_input_bits_31; // @[TCU.scala 71:19]
  wire  mem_io_portA_output_ready; // @[TCU.scala 71:19]
  wire  mem_io_portA_output_valid; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_0; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_1; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_2; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_3; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_4; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_5; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_6; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_7; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_8; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_9; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_10; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_11; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_12; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_13; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_14; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_15; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_16; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_17; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_18; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_19; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_20; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_21; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_22; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_23; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_24; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_25; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_26; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_27; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_28; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_29; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_30; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portA_output_bits_31; // @[TCU.scala 71:19]
  wire  mem_io_portB_control_ready; // @[TCU.scala 71:19]
  wire  mem_io_portB_control_valid; // @[TCU.scala 71:19]
  wire  mem_io_portB_control_bits_write; // @[TCU.scala 71:19]
  wire [13:0] mem_io_portB_control_bits_address; // @[TCU.scala 71:19]
  wire  mem_io_portB_input_ready; // @[TCU.scala 71:19]
  wire  mem_io_portB_input_valid; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_0; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_1; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_2; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_3; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_4; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_5; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_6; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_7; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_8; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_9; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_10; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_11; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_12; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_13; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_14; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_15; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_16; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_17; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_18; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_19; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_20; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_21; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_22; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_23; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_24; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_25; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_26; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_27; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_28; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_29; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_30; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_input_bits_31; // @[TCU.scala 71:19]
  wire  mem_io_portB_output_ready; // @[TCU.scala 71:19]
  wire  mem_io_portB_output_valid; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_0; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_1; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_2; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_3; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_4; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_5; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_6; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_7; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_8; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_9; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_10; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_11; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_12; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_13; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_14; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_15; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_16; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_17; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_18; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_19; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_20; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_21; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_22; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_23; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_24; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_25; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_26; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_27; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_28; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_29; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_30; // @[TCU.scala 71:19]
  wire [15:0] mem_io_portB_output_bits_31; // @[TCU.scala 71:19]
  wire  mem_io_tracepoint; // @[TCU.scala 71:19]
  wire [31:0] mem_io_programCounter; // @[TCU.scala 71:19]
  wire  router_clock; // @[TCU.scala 80:22]
  wire  router_reset; // @[TCU.scala 80:22]
  wire  router_io_control_ready; // @[TCU.scala 80:22]
  wire  router_io_control_valid; // @[TCU.scala 80:22]
  wire [3:0] router_io_control_bits_kind; // @[TCU.scala 80:22]
  wire [13:0] router_io_control_bits_size; // @[TCU.scala 80:22]
  wire  router_io_mem_output_ready; // @[TCU.scala 80:22]
  wire  router_io_mem_output_valid; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_0; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_1; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_2; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_3; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_4; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_5; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_6; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_7; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_8; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_9; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_10; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_11; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_12; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_13; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_14; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_15; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_16; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_17; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_18; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_19; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_20; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_21; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_22; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_23; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_24; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_25; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_26; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_27; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_28; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_29; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_30; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_output_bits_31; // @[TCU.scala 80:22]
  wire  router_io_mem_input_ready; // @[TCU.scala 80:22]
  wire  router_io_mem_input_valid; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_0; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_1; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_2; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_3; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_4; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_5; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_6; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_7; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_8; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_9; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_10; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_11; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_12; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_13; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_14; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_15; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_16; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_17; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_18; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_19; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_20; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_21; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_22; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_23; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_24; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_25; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_26; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_27; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_28; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_29; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_30; // @[TCU.scala 80:22]
  wire [15:0] router_io_mem_input_bits_31; // @[TCU.scala 80:22]
  wire  router_io_array_input_ready; // @[TCU.scala 80:22]
  wire  router_io_array_input_valid; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_0; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_1; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_2; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_3; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_4; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_5; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_6; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_7; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_8; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_9; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_10; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_11; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_12; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_13; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_14; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_15; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_16; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_17; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_18; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_19; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_20; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_21; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_22; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_23; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_24; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_25; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_26; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_27; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_28; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_29; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_30; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_input_bits_31; // @[TCU.scala 80:22]
  wire  router_io_array_output_ready; // @[TCU.scala 80:22]
  wire  router_io_array_output_valid; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_0; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_1; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_2; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_3; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_4; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_5; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_6; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_7; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_8; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_9; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_10; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_11; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_12; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_13; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_14; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_15; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_16; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_17; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_18; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_19; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_20; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_21; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_22; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_23; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_24; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_25; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_26; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_27; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_28; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_29; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_30; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_output_bits_31; // @[TCU.scala 80:22]
  wire  router_io_array_weightInput_ready; // @[TCU.scala 80:22]
  wire  router_io_array_weightInput_valid; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_0; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_1; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_2; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_3; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_4; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_5; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_6; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_7; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_8; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_9; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_10; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_11; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_12; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_13; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_14; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_15; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_16; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_17; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_18; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_19; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_20; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_21; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_22; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_23; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_24; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_25; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_26; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_27; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_28; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_29; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_30; // @[TCU.scala 80:22]
  wire [15:0] router_io_array_weightInput_bits_31; // @[TCU.scala 80:22]
  wire  router_io_acc_output_ready; // @[TCU.scala 80:22]
  wire  router_io_acc_output_valid; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_0; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_1; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_2; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_3; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_4; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_5; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_6; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_7; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_8; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_9; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_10; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_11; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_12; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_13; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_14; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_15; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_16; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_17; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_18; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_19; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_20; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_21; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_22; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_23; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_24; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_25; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_26; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_27; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_28; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_29; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_30; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_output_bits_31; // @[TCU.scala 80:22]
  wire  router_io_acc_input_ready; // @[TCU.scala 80:22]
  wire  router_io_acc_input_valid; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_0; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_1; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_2; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_3; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_4; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_5; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_6; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_7; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_8; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_9; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_10; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_11; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_12; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_13; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_14; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_15; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_16; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_17; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_18; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_19; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_20; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_21; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_22; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_23; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_24; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_25; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_26; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_27; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_28; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_29; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_30; // @[TCU.scala 80:22]
  wire [15:0] router_io_acc_input_bits_31; // @[TCU.scala 80:22]
  wire  router_io_timeout; // @[TCU.scala 80:22]
  wire  router_io_tracepoint; // @[TCU.scala 80:22]
  wire [31:0] router_io_programCounter; // @[TCU.scala 80:22]
  wire  hostRouter_io_control_ready; // @[TCU.scala 87:26]
  wire  hostRouter_io_control_valid; // @[TCU.scala 87:26]
  wire [1:0] hostRouter_io_control_bits_kind; // @[TCU.scala 87:26]
  wire  hostRouter_io_dram0_dataIn_ready; // @[TCU.scala 87:26]
  wire  hostRouter_io_dram0_dataIn_valid; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_0; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_1; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_2; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_3; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_4; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_5; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_6; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_7; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_8; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_9; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_10; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_11; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_12; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_13; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_14; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_15; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_16; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_17; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_18; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_19; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_20; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_21; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_22; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_23; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_24; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_25; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_26; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_27; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_28; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_29; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_30; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataIn_bits_31; // @[TCU.scala 87:26]
  wire  hostRouter_io_dram0_dataOut_ready; // @[TCU.scala 87:26]
  wire  hostRouter_io_dram0_dataOut_valid; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_0; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_1; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_2; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_3; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_4; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_5; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_6; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_7; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_8; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_9; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_10; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_11; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_12; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_13; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_14; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_15; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_16; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_17; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_18; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_19; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_20; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_21; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_22; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_23; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_24; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_25; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_26; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_27; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_28; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_29; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_30; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram0_dataOut_bits_31; // @[TCU.scala 87:26]
  wire  hostRouter_io_dram1_dataIn_ready; // @[TCU.scala 87:26]
  wire  hostRouter_io_dram1_dataIn_valid; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_0; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_1; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_2; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_3; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_4; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_5; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_6; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_7; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_8; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_9; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_10; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_11; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_12; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_13; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_14; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_15; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_16; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_17; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_18; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_19; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_20; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_21; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_22; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_23; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_24; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_25; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_26; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_27; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_28; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_29; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_30; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataIn_bits_31; // @[TCU.scala 87:26]
  wire  hostRouter_io_dram1_dataOut_ready; // @[TCU.scala 87:26]
  wire  hostRouter_io_dram1_dataOut_valid; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_0; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_1; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_2; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_3; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_4; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_5; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_6; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_7; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_8; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_9; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_10; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_11; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_12; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_13; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_14; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_15; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_16; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_17; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_18; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_19; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_20; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_21; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_22; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_23; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_24; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_25; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_26; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_27; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_28; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_29; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_30; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_dram1_dataOut_bits_31; // @[TCU.scala 87:26]
  wire  hostRouter_io_mem_output_ready; // @[TCU.scala 87:26]
  wire  hostRouter_io_mem_output_valid; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_0; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_1; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_2; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_3; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_4; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_5; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_6; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_7; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_8; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_9; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_10; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_11; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_12; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_13; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_14; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_15; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_16; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_17; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_18; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_19; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_20; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_21; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_22; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_23; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_24; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_25; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_26; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_27; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_28; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_29; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_30; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_output_bits_31; // @[TCU.scala 87:26]
  wire  hostRouter_io_mem_input_ready; // @[TCU.scala 87:26]
  wire  hostRouter_io_mem_input_valid; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_0; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_1; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_2; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_3; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_4; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_5; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_6; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_7; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_8; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_9; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_10; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_11; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_12; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_13; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_14; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_15; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_16; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_17; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_18; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_19; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_20; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_21; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_22; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_23; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_24; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_25; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_26; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_27; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_28; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_29; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_30; // @[TCU.scala 87:26]
  wire [15:0] hostRouter_io_mem_input_bits_31; // @[TCU.scala 87:26]
  wire  acc_io_control_q_clock; // @[TCU.scala 110:39]
  wire  acc_io_control_q_reset; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_enq_ready; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_enq_valid; // @[TCU.scala 110:39]
  wire [3:0] acc_io_control_q_io_enq_bits_instruction_op; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_enq_bits_instruction_sourceLeft; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_enq_bits_instruction_sourceRight; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_enq_bits_instruction_dest; // @[TCU.scala 110:39]
  wire [11:0] acc_io_control_q_io_enq_bits_readAddress; // @[TCU.scala 110:39]
  wire [11:0] acc_io_control_q_io_enq_bits_writeAddress; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_enq_bits_accumulate; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_enq_bits_write; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_enq_bits_read; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_deq_ready; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_deq_valid; // @[TCU.scala 110:39]
  wire [3:0] acc_io_control_q_io_deq_bits_instruction_op; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_deq_bits_instruction_sourceLeft; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_deq_bits_instruction_sourceRight; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_deq_bits_instruction_dest; // @[TCU.scala 110:39]
  wire [11:0] acc_io_control_q_io_deq_bits_readAddress; // @[TCU.scala 110:39]
  wire [11:0] acc_io_control_q_io_deq_bits_writeAddress; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_deq_bits_accumulate; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_deq_bits_write; // @[TCU.scala 110:39]
  wire  acc_io_control_q_io_deq_bits_read; // @[TCU.scala 110:39]
  wire  array_io_control_q_clock; // @[TCU.scala 117:41]
  wire  array_io_control_q_reset; // @[TCU.scala 117:41]
  wire  array_io_control_q_io_enq_ready; // @[TCU.scala 117:41]
  wire  array_io_control_q_io_enq_valid; // @[TCU.scala 117:41]
  wire  array_io_control_q_io_enq_bits_load; // @[TCU.scala 117:41]
  wire  array_io_control_q_io_enq_bits_zeroes; // @[TCU.scala 117:41]
  wire  array_io_control_q_io_deq_ready; // @[TCU.scala 117:41]
  wire  array_io_control_q_io_deq_valid; // @[TCU.scala 117:41]
  wire  array_io_control_q_io_deq_bits_load; // @[TCU.scala 117:41]
  wire  array_io_control_q_io_deq_bits_zeroes; // @[TCU.scala 117:41]
  Decoder decoder ( // @[TCU.scala 64:23]
    .clock(decoder_clock),
    .reset(decoder_reset),
    .io_instruction_ready(decoder_io_instruction_ready),
    .io_instruction_valid(decoder_io_instruction_valid),
    .io_instruction_bits_opcode(decoder_io_instruction_bits_opcode),
    .io_instruction_bits_flags(decoder_io_instruction_bits_flags),
    .io_instruction_bits_arguments(decoder_io_instruction_bits_arguments),
    .io_memPortA_ready(decoder_io_memPortA_ready),
    .io_memPortA_valid(decoder_io_memPortA_valid),
    .io_memPortA_bits_write(decoder_io_memPortA_bits_write),
    .io_memPortA_bits_address(decoder_io_memPortA_bits_address),
    .io_memPortB_ready(decoder_io_memPortB_ready),
    .io_memPortB_valid(decoder_io_memPortB_valid),
    .io_memPortB_bits_write(decoder_io_memPortB_bits_write),
    .io_memPortB_bits_address(decoder_io_memPortB_bits_address),
    .io_dram0_ready(decoder_io_dram0_ready),
    .io_dram0_valid(decoder_io_dram0_valid),
    .io_dram0_bits_write(decoder_io_dram0_bits_write),
    .io_dram0_bits_address(decoder_io_dram0_bits_address),
    .io_dram0_bits_size(decoder_io_dram0_bits_size),
    .io_dram1_ready(decoder_io_dram1_ready),
    .io_dram1_valid(decoder_io_dram1_valid),
    .io_dram1_bits_write(decoder_io_dram1_bits_write),
    .io_dram1_bits_address(decoder_io_dram1_bits_address),
    .io_dram1_bits_size(decoder_io_dram1_bits_size),
    .io_dataflow_ready(decoder_io_dataflow_ready),
    .io_dataflow_valid(decoder_io_dataflow_valid),
    .io_dataflow_bits_kind(decoder_io_dataflow_bits_kind),
    .io_dataflow_bits_size(decoder_io_dataflow_bits_size),
    .io_hostDataflow_ready(decoder_io_hostDataflow_ready),
    .io_hostDataflow_valid(decoder_io_hostDataflow_valid),
    .io_hostDataflow_bits_kind(decoder_io_hostDataflow_bits_kind),
    .io_acc_ready(decoder_io_acc_ready),
    .io_acc_valid(decoder_io_acc_valid),
    .io_acc_bits_instruction_op(decoder_io_acc_bits_instruction_op),
    .io_acc_bits_instruction_sourceLeft(decoder_io_acc_bits_instruction_sourceLeft),
    .io_acc_bits_instruction_sourceRight(decoder_io_acc_bits_instruction_sourceRight),
    .io_acc_bits_instruction_dest(decoder_io_acc_bits_instruction_dest),
    .io_acc_bits_readAddress(decoder_io_acc_bits_readAddress),
    .io_acc_bits_writeAddress(decoder_io_acc_bits_writeAddress),
    .io_acc_bits_accumulate(decoder_io_acc_bits_accumulate),
    .io_acc_bits_write(decoder_io_acc_bits_write),
    .io_acc_bits_read(decoder_io_acc_bits_read),
    .io_array_ready(decoder_io_array_ready),
    .io_array_valid(decoder_io_array_valid),
    .io_array_bits_load(decoder_io_array_bits_load),
    .io_array_bits_zeroes(decoder_io_array_bits_zeroes),
    .io_config_dram0AddressOffset(decoder_io_config_dram0AddressOffset),
    .io_config_dram0CacheBehaviour(decoder_io_config_dram0CacheBehaviour),
    .io_config_dram1AddressOffset(decoder_io_config_dram1AddressOffset),
    .io_config_dram1CacheBehaviour(decoder_io_config_dram1CacheBehaviour),
    .io_timeout(decoder_io_timeout),
    .io_error(decoder_io_error),
    .io_tracepoint(decoder_io_tracepoint),
    .io_programCounter(decoder_io_programCounter)
  );
  SystolicArray array ( // @[TCU.scala 65:21]
    .clock(array_clock),
    .reset(array_reset),
    .io_control_ready(array_io_control_ready),
    .io_control_valid(array_io_control_valid),
    .io_control_bits_load(array_io_control_bits_load),
    .io_control_bits_zeroes(array_io_control_bits_zeroes),
    .io_input_ready(array_io_input_ready),
    .io_input_valid(array_io_input_valid),
    .io_input_bits_0(array_io_input_bits_0),
    .io_input_bits_1(array_io_input_bits_1),
    .io_input_bits_2(array_io_input_bits_2),
    .io_input_bits_3(array_io_input_bits_3),
    .io_input_bits_4(array_io_input_bits_4),
    .io_input_bits_5(array_io_input_bits_5),
    .io_input_bits_6(array_io_input_bits_6),
    .io_input_bits_7(array_io_input_bits_7),
    .io_input_bits_8(array_io_input_bits_8),
    .io_input_bits_9(array_io_input_bits_9),
    .io_input_bits_10(array_io_input_bits_10),
    .io_input_bits_11(array_io_input_bits_11),
    .io_input_bits_12(array_io_input_bits_12),
    .io_input_bits_13(array_io_input_bits_13),
    .io_input_bits_14(array_io_input_bits_14),
    .io_input_bits_15(array_io_input_bits_15),
    .io_input_bits_16(array_io_input_bits_16),
    .io_input_bits_17(array_io_input_bits_17),
    .io_input_bits_18(array_io_input_bits_18),
    .io_input_bits_19(array_io_input_bits_19),
    .io_input_bits_20(array_io_input_bits_20),
    .io_input_bits_21(array_io_input_bits_21),
    .io_input_bits_22(array_io_input_bits_22),
    .io_input_bits_23(array_io_input_bits_23),
    .io_input_bits_24(array_io_input_bits_24),
    .io_input_bits_25(array_io_input_bits_25),
    .io_input_bits_26(array_io_input_bits_26),
    .io_input_bits_27(array_io_input_bits_27),
    .io_input_bits_28(array_io_input_bits_28),
    .io_input_bits_29(array_io_input_bits_29),
    .io_input_bits_30(array_io_input_bits_30),
    .io_input_bits_31(array_io_input_bits_31),
    .io_weight_ready(array_io_weight_ready),
    .io_weight_valid(array_io_weight_valid),
    .io_weight_bits_0(array_io_weight_bits_0),
    .io_weight_bits_1(array_io_weight_bits_1),
    .io_weight_bits_2(array_io_weight_bits_2),
    .io_weight_bits_3(array_io_weight_bits_3),
    .io_weight_bits_4(array_io_weight_bits_4),
    .io_weight_bits_5(array_io_weight_bits_5),
    .io_weight_bits_6(array_io_weight_bits_6),
    .io_weight_bits_7(array_io_weight_bits_7),
    .io_weight_bits_8(array_io_weight_bits_8),
    .io_weight_bits_9(array_io_weight_bits_9),
    .io_weight_bits_10(array_io_weight_bits_10),
    .io_weight_bits_11(array_io_weight_bits_11),
    .io_weight_bits_12(array_io_weight_bits_12),
    .io_weight_bits_13(array_io_weight_bits_13),
    .io_weight_bits_14(array_io_weight_bits_14),
    .io_weight_bits_15(array_io_weight_bits_15),
    .io_weight_bits_16(array_io_weight_bits_16),
    .io_weight_bits_17(array_io_weight_bits_17),
    .io_weight_bits_18(array_io_weight_bits_18),
    .io_weight_bits_19(array_io_weight_bits_19),
    .io_weight_bits_20(array_io_weight_bits_20),
    .io_weight_bits_21(array_io_weight_bits_21),
    .io_weight_bits_22(array_io_weight_bits_22),
    .io_weight_bits_23(array_io_weight_bits_23),
    .io_weight_bits_24(array_io_weight_bits_24),
    .io_weight_bits_25(array_io_weight_bits_25),
    .io_weight_bits_26(array_io_weight_bits_26),
    .io_weight_bits_27(array_io_weight_bits_27),
    .io_weight_bits_28(array_io_weight_bits_28),
    .io_weight_bits_29(array_io_weight_bits_29),
    .io_weight_bits_30(array_io_weight_bits_30),
    .io_weight_bits_31(array_io_weight_bits_31),
    .io_output_ready(array_io_output_ready),
    .io_output_valid(array_io_output_valid),
    .io_output_bits_0(array_io_output_bits_0),
    .io_output_bits_1(array_io_output_bits_1),
    .io_output_bits_2(array_io_output_bits_2),
    .io_output_bits_3(array_io_output_bits_3),
    .io_output_bits_4(array_io_output_bits_4),
    .io_output_bits_5(array_io_output_bits_5),
    .io_output_bits_6(array_io_output_bits_6),
    .io_output_bits_7(array_io_output_bits_7),
    .io_output_bits_8(array_io_output_bits_8),
    .io_output_bits_9(array_io_output_bits_9),
    .io_output_bits_10(array_io_output_bits_10),
    .io_output_bits_11(array_io_output_bits_11),
    .io_output_bits_12(array_io_output_bits_12),
    .io_output_bits_13(array_io_output_bits_13),
    .io_output_bits_14(array_io_output_bits_14),
    .io_output_bits_15(array_io_output_bits_15),
    .io_output_bits_16(array_io_output_bits_16),
    .io_output_bits_17(array_io_output_bits_17),
    .io_output_bits_18(array_io_output_bits_18),
    .io_output_bits_19(array_io_output_bits_19),
    .io_output_bits_20(array_io_output_bits_20),
    .io_output_bits_21(array_io_output_bits_21),
    .io_output_bits_22(array_io_output_bits_22),
    .io_output_bits_23(array_io_output_bits_23),
    .io_output_bits_24(array_io_output_bits_24),
    .io_output_bits_25(array_io_output_bits_25),
    .io_output_bits_26(array_io_output_bits_26),
    .io_output_bits_27(array_io_output_bits_27),
    .io_output_bits_28(array_io_output_bits_28),
    .io_output_bits_29(array_io_output_bits_29),
    .io_output_bits_30(array_io_output_bits_30),
    .io_output_bits_31(array_io_output_bits_31)
  );
  AccumulatorWithALUArray acc ( // @[TCU.scala 68:19]
    .clock(acc_clock),
    .reset(acc_reset),
    .io_input_ready(acc_io_input_ready),
    .io_input_valid(acc_io_input_valid),
    .io_input_bits_0(acc_io_input_bits_0),
    .io_input_bits_1(acc_io_input_bits_1),
    .io_input_bits_2(acc_io_input_bits_2),
    .io_input_bits_3(acc_io_input_bits_3),
    .io_input_bits_4(acc_io_input_bits_4),
    .io_input_bits_5(acc_io_input_bits_5),
    .io_input_bits_6(acc_io_input_bits_6),
    .io_input_bits_7(acc_io_input_bits_7),
    .io_input_bits_8(acc_io_input_bits_8),
    .io_input_bits_9(acc_io_input_bits_9),
    .io_input_bits_10(acc_io_input_bits_10),
    .io_input_bits_11(acc_io_input_bits_11),
    .io_input_bits_12(acc_io_input_bits_12),
    .io_input_bits_13(acc_io_input_bits_13),
    .io_input_bits_14(acc_io_input_bits_14),
    .io_input_bits_15(acc_io_input_bits_15),
    .io_input_bits_16(acc_io_input_bits_16),
    .io_input_bits_17(acc_io_input_bits_17),
    .io_input_bits_18(acc_io_input_bits_18),
    .io_input_bits_19(acc_io_input_bits_19),
    .io_input_bits_20(acc_io_input_bits_20),
    .io_input_bits_21(acc_io_input_bits_21),
    .io_input_bits_22(acc_io_input_bits_22),
    .io_input_bits_23(acc_io_input_bits_23),
    .io_input_bits_24(acc_io_input_bits_24),
    .io_input_bits_25(acc_io_input_bits_25),
    .io_input_bits_26(acc_io_input_bits_26),
    .io_input_bits_27(acc_io_input_bits_27),
    .io_input_bits_28(acc_io_input_bits_28),
    .io_input_bits_29(acc_io_input_bits_29),
    .io_input_bits_30(acc_io_input_bits_30),
    .io_input_bits_31(acc_io_input_bits_31),
    .io_output_ready(acc_io_output_ready),
    .io_output_valid(acc_io_output_valid),
    .io_output_bits_0(acc_io_output_bits_0),
    .io_output_bits_1(acc_io_output_bits_1),
    .io_output_bits_2(acc_io_output_bits_2),
    .io_output_bits_3(acc_io_output_bits_3),
    .io_output_bits_4(acc_io_output_bits_4),
    .io_output_bits_5(acc_io_output_bits_5),
    .io_output_bits_6(acc_io_output_bits_6),
    .io_output_bits_7(acc_io_output_bits_7),
    .io_output_bits_8(acc_io_output_bits_8),
    .io_output_bits_9(acc_io_output_bits_9),
    .io_output_bits_10(acc_io_output_bits_10),
    .io_output_bits_11(acc_io_output_bits_11),
    .io_output_bits_12(acc_io_output_bits_12),
    .io_output_bits_13(acc_io_output_bits_13),
    .io_output_bits_14(acc_io_output_bits_14),
    .io_output_bits_15(acc_io_output_bits_15),
    .io_output_bits_16(acc_io_output_bits_16),
    .io_output_bits_17(acc_io_output_bits_17),
    .io_output_bits_18(acc_io_output_bits_18),
    .io_output_bits_19(acc_io_output_bits_19),
    .io_output_bits_20(acc_io_output_bits_20),
    .io_output_bits_21(acc_io_output_bits_21),
    .io_output_bits_22(acc_io_output_bits_22),
    .io_output_bits_23(acc_io_output_bits_23),
    .io_output_bits_24(acc_io_output_bits_24),
    .io_output_bits_25(acc_io_output_bits_25),
    .io_output_bits_26(acc_io_output_bits_26),
    .io_output_bits_27(acc_io_output_bits_27),
    .io_output_bits_28(acc_io_output_bits_28),
    .io_output_bits_29(acc_io_output_bits_29),
    .io_output_bits_30(acc_io_output_bits_30),
    .io_output_bits_31(acc_io_output_bits_31),
    .io_control_ready(acc_io_control_ready),
    .io_control_valid(acc_io_control_valid),
    .io_control_bits_instruction_op(acc_io_control_bits_instruction_op),
    .io_control_bits_instruction_sourceLeft(acc_io_control_bits_instruction_sourceLeft),
    .io_control_bits_instruction_sourceRight(acc_io_control_bits_instruction_sourceRight),
    .io_control_bits_instruction_dest(acc_io_control_bits_instruction_dest),
    .io_control_bits_readAddress(acc_io_control_bits_readAddress),
    .io_control_bits_writeAddress(acc_io_control_bits_writeAddress),
    .io_control_bits_accumulate(acc_io_control_bits_accumulate),
    .io_control_bits_write(acc_io_control_bits_write),
    .io_control_bits_read(acc_io_control_bits_read),
    .io_tracepoint(acc_io_tracepoint),
    .io_programCounter(acc_io_programCounter)
  );
  DualPortMem_1 mem ( // @[TCU.scala 71:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_portA_control_ready(mem_io_portA_control_ready),
    .io_portA_control_valid(mem_io_portA_control_valid),
    .io_portA_control_bits_write(mem_io_portA_control_bits_write),
    .io_portA_control_bits_address(mem_io_portA_control_bits_address),
    .io_portA_input_ready(mem_io_portA_input_ready),
    .io_portA_input_valid(mem_io_portA_input_valid),
    .io_portA_input_bits_0(mem_io_portA_input_bits_0),
    .io_portA_input_bits_1(mem_io_portA_input_bits_1),
    .io_portA_input_bits_2(mem_io_portA_input_bits_2),
    .io_portA_input_bits_3(mem_io_portA_input_bits_3),
    .io_portA_input_bits_4(mem_io_portA_input_bits_4),
    .io_portA_input_bits_5(mem_io_portA_input_bits_5),
    .io_portA_input_bits_6(mem_io_portA_input_bits_6),
    .io_portA_input_bits_7(mem_io_portA_input_bits_7),
    .io_portA_input_bits_8(mem_io_portA_input_bits_8),
    .io_portA_input_bits_9(mem_io_portA_input_bits_9),
    .io_portA_input_bits_10(mem_io_portA_input_bits_10),
    .io_portA_input_bits_11(mem_io_portA_input_bits_11),
    .io_portA_input_bits_12(mem_io_portA_input_bits_12),
    .io_portA_input_bits_13(mem_io_portA_input_bits_13),
    .io_portA_input_bits_14(mem_io_portA_input_bits_14),
    .io_portA_input_bits_15(mem_io_portA_input_bits_15),
    .io_portA_input_bits_16(mem_io_portA_input_bits_16),
    .io_portA_input_bits_17(mem_io_portA_input_bits_17),
    .io_portA_input_bits_18(mem_io_portA_input_bits_18),
    .io_portA_input_bits_19(mem_io_portA_input_bits_19),
    .io_portA_input_bits_20(mem_io_portA_input_bits_20),
    .io_portA_input_bits_21(mem_io_portA_input_bits_21),
    .io_portA_input_bits_22(mem_io_portA_input_bits_22),
    .io_portA_input_bits_23(mem_io_portA_input_bits_23),
    .io_portA_input_bits_24(mem_io_portA_input_bits_24),
    .io_portA_input_bits_25(mem_io_portA_input_bits_25),
    .io_portA_input_bits_26(mem_io_portA_input_bits_26),
    .io_portA_input_bits_27(mem_io_portA_input_bits_27),
    .io_portA_input_bits_28(mem_io_portA_input_bits_28),
    .io_portA_input_bits_29(mem_io_portA_input_bits_29),
    .io_portA_input_bits_30(mem_io_portA_input_bits_30),
    .io_portA_input_bits_31(mem_io_portA_input_bits_31),
    .io_portA_output_ready(mem_io_portA_output_ready),
    .io_portA_output_valid(mem_io_portA_output_valid),
    .io_portA_output_bits_0(mem_io_portA_output_bits_0),
    .io_portA_output_bits_1(mem_io_portA_output_bits_1),
    .io_portA_output_bits_2(mem_io_portA_output_bits_2),
    .io_portA_output_bits_3(mem_io_portA_output_bits_3),
    .io_portA_output_bits_4(mem_io_portA_output_bits_4),
    .io_portA_output_bits_5(mem_io_portA_output_bits_5),
    .io_portA_output_bits_6(mem_io_portA_output_bits_6),
    .io_portA_output_bits_7(mem_io_portA_output_bits_7),
    .io_portA_output_bits_8(mem_io_portA_output_bits_8),
    .io_portA_output_bits_9(mem_io_portA_output_bits_9),
    .io_portA_output_bits_10(mem_io_portA_output_bits_10),
    .io_portA_output_bits_11(mem_io_portA_output_bits_11),
    .io_portA_output_bits_12(mem_io_portA_output_bits_12),
    .io_portA_output_bits_13(mem_io_portA_output_bits_13),
    .io_portA_output_bits_14(mem_io_portA_output_bits_14),
    .io_portA_output_bits_15(mem_io_portA_output_bits_15),
    .io_portA_output_bits_16(mem_io_portA_output_bits_16),
    .io_portA_output_bits_17(mem_io_portA_output_bits_17),
    .io_portA_output_bits_18(mem_io_portA_output_bits_18),
    .io_portA_output_bits_19(mem_io_portA_output_bits_19),
    .io_portA_output_bits_20(mem_io_portA_output_bits_20),
    .io_portA_output_bits_21(mem_io_portA_output_bits_21),
    .io_portA_output_bits_22(mem_io_portA_output_bits_22),
    .io_portA_output_bits_23(mem_io_portA_output_bits_23),
    .io_portA_output_bits_24(mem_io_portA_output_bits_24),
    .io_portA_output_bits_25(mem_io_portA_output_bits_25),
    .io_portA_output_bits_26(mem_io_portA_output_bits_26),
    .io_portA_output_bits_27(mem_io_portA_output_bits_27),
    .io_portA_output_bits_28(mem_io_portA_output_bits_28),
    .io_portA_output_bits_29(mem_io_portA_output_bits_29),
    .io_portA_output_bits_30(mem_io_portA_output_bits_30),
    .io_portA_output_bits_31(mem_io_portA_output_bits_31),
    .io_portB_control_ready(mem_io_portB_control_ready),
    .io_portB_control_valid(mem_io_portB_control_valid),
    .io_portB_control_bits_write(mem_io_portB_control_bits_write),
    .io_portB_control_bits_address(mem_io_portB_control_bits_address),
    .io_portB_input_ready(mem_io_portB_input_ready),
    .io_portB_input_valid(mem_io_portB_input_valid),
    .io_portB_input_bits_0(mem_io_portB_input_bits_0),
    .io_portB_input_bits_1(mem_io_portB_input_bits_1),
    .io_portB_input_bits_2(mem_io_portB_input_bits_2),
    .io_portB_input_bits_3(mem_io_portB_input_bits_3),
    .io_portB_input_bits_4(mem_io_portB_input_bits_4),
    .io_portB_input_bits_5(mem_io_portB_input_bits_5),
    .io_portB_input_bits_6(mem_io_portB_input_bits_6),
    .io_portB_input_bits_7(mem_io_portB_input_bits_7),
    .io_portB_input_bits_8(mem_io_portB_input_bits_8),
    .io_portB_input_bits_9(mem_io_portB_input_bits_9),
    .io_portB_input_bits_10(mem_io_portB_input_bits_10),
    .io_portB_input_bits_11(mem_io_portB_input_bits_11),
    .io_portB_input_bits_12(mem_io_portB_input_bits_12),
    .io_portB_input_bits_13(mem_io_portB_input_bits_13),
    .io_portB_input_bits_14(mem_io_portB_input_bits_14),
    .io_portB_input_bits_15(mem_io_portB_input_bits_15),
    .io_portB_input_bits_16(mem_io_portB_input_bits_16),
    .io_portB_input_bits_17(mem_io_portB_input_bits_17),
    .io_portB_input_bits_18(mem_io_portB_input_bits_18),
    .io_portB_input_bits_19(mem_io_portB_input_bits_19),
    .io_portB_input_bits_20(mem_io_portB_input_bits_20),
    .io_portB_input_bits_21(mem_io_portB_input_bits_21),
    .io_portB_input_bits_22(mem_io_portB_input_bits_22),
    .io_portB_input_bits_23(mem_io_portB_input_bits_23),
    .io_portB_input_bits_24(mem_io_portB_input_bits_24),
    .io_portB_input_bits_25(mem_io_portB_input_bits_25),
    .io_portB_input_bits_26(mem_io_portB_input_bits_26),
    .io_portB_input_bits_27(mem_io_portB_input_bits_27),
    .io_portB_input_bits_28(mem_io_portB_input_bits_28),
    .io_portB_input_bits_29(mem_io_portB_input_bits_29),
    .io_portB_input_bits_30(mem_io_portB_input_bits_30),
    .io_portB_input_bits_31(mem_io_portB_input_bits_31),
    .io_portB_output_ready(mem_io_portB_output_ready),
    .io_portB_output_valid(mem_io_portB_output_valid),
    .io_portB_output_bits_0(mem_io_portB_output_bits_0),
    .io_portB_output_bits_1(mem_io_portB_output_bits_1),
    .io_portB_output_bits_2(mem_io_portB_output_bits_2),
    .io_portB_output_bits_3(mem_io_portB_output_bits_3),
    .io_portB_output_bits_4(mem_io_portB_output_bits_4),
    .io_portB_output_bits_5(mem_io_portB_output_bits_5),
    .io_portB_output_bits_6(mem_io_portB_output_bits_6),
    .io_portB_output_bits_7(mem_io_portB_output_bits_7),
    .io_portB_output_bits_8(mem_io_portB_output_bits_8),
    .io_portB_output_bits_9(mem_io_portB_output_bits_9),
    .io_portB_output_bits_10(mem_io_portB_output_bits_10),
    .io_portB_output_bits_11(mem_io_portB_output_bits_11),
    .io_portB_output_bits_12(mem_io_portB_output_bits_12),
    .io_portB_output_bits_13(mem_io_portB_output_bits_13),
    .io_portB_output_bits_14(mem_io_portB_output_bits_14),
    .io_portB_output_bits_15(mem_io_portB_output_bits_15),
    .io_portB_output_bits_16(mem_io_portB_output_bits_16),
    .io_portB_output_bits_17(mem_io_portB_output_bits_17),
    .io_portB_output_bits_18(mem_io_portB_output_bits_18),
    .io_portB_output_bits_19(mem_io_portB_output_bits_19),
    .io_portB_output_bits_20(mem_io_portB_output_bits_20),
    .io_portB_output_bits_21(mem_io_portB_output_bits_21),
    .io_portB_output_bits_22(mem_io_portB_output_bits_22),
    .io_portB_output_bits_23(mem_io_portB_output_bits_23),
    .io_portB_output_bits_24(mem_io_portB_output_bits_24),
    .io_portB_output_bits_25(mem_io_portB_output_bits_25),
    .io_portB_output_bits_26(mem_io_portB_output_bits_26),
    .io_portB_output_bits_27(mem_io_portB_output_bits_27),
    .io_portB_output_bits_28(mem_io_portB_output_bits_28),
    .io_portB_output_bits_29(mem_io_portB_output_bits_29),
    .io_portB_output_bits_30(mem_io_portB_output_bits_30),
    .io_portB_output_bits_31(mem_io_portB_output_bits_31),
    .io_tracepoint(mem_io_tracepoint),
    .io_programCounter(mem_io_programCounter)
  );
  LocalRouter router ( // @[TCU.scala 80:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_control_ready(router_io_control_ready),
    .io_control_valid(router_io_control_valid),
    .io_control_bits_kind(router_io_control_bits_kind),
    .io_control_bits_size(router_io_control_bits_size),
    .io_mem_output_ready(router_io_mem_output_ready),
    .io_mem_output_valid(router_io_mem_output_valid),
    .io_mem_output_bits_0(router_io_mem_output_bits_0),
    .io_mem_output_bits_1(router_io_mem_output_bits_1),
    .io_mem_output_bits_2(router_io_mem_output_bits_2),
    .io_mem_output_bits_3(router_io_mem_output_bits_3),
    .io_mem_output_bits_4(router_io_mem_output_bits_4),
    .io_mem_output_bits_5(router_io_mem_output_bits_5),
    .io_mem_output_bits_6(router_io_mem_output_bits_6),
    .io_mem_output_bits_7(router_io_mem_output_bits_7),
    .io_mem_output_bits_8(router_io_mem_output_bits_8),
    .io_mem_output_bits_9(router_io_mem_output_bits_9),
    .io_mem_output_bits_10(router_io_mem_output_bits_10),
    .io_mem_output_bits_11(router_io_mem_output_bits_11),
    .io_mem_output_bits_12(router_io_mem_output_bits_12),
    .io_mem_output_bits_13(router_io_mem_output_bits_13),
    .io_mem_output_bits_14(router_io_mem_output_bits_14),
    .io_mem_output_bits_15(router_io_mem_output_bits_15),
    .io_mem_output_bits_16(router_io_mem_output_bits_16),
    .io_mem_output_bits_17(router_io_mem_output_bits_17),
    .io_mem_output_bits_18(router_io_mem_output_bits_18),
    .io_mem_output_bits_19(router_io_mem_output_bits_19),
    .io_mem_output_bits_20(router_io_mem_output_bits_20),
    .io_mem_output_bits_21(router_io_mem_output_bits_21),
    .io_mem_output_bits_22(router_io_mem_output_bits_22),
    .io_mem_output_bits_23(router_io_mem_output_bits_23),
    .io_mem_output_bits_24(router_io_mem_output_bits_24),
    .io_mem_output_bits_25(router_io_mem_output_bits_25),
    .io_mem_output_bits_26(router_io_mem_output_bits_26),
    .io_mem_output_bits_27(router_io_mem_output_bits_27),
    .io_mem_output_bits_28(router_io_mem_output_bits_28),
    .io_mem_output_bits_29(router_io_mem_output_bits_29),
    .io_mem_output_bits_30(router_io_mem_output_bits_30),
    .io_mem_output_bits_31(router_io_mem_output_bits_31),
    .io_mem_input_ready(router_io_mem_input_ready),
    .io_mem_input_valid(router_io_mem_input_valid),
    .io_mem_input_bits_0(router_io_mem_input_bits_0),
    .io_mem_input_bits_1(router_io_mem_input_bits_1),
    .io_mem_input_bits_2(router_io_mem_input_bits_2),
    .io_mem_input_bits_3(router_io_mem_input_bits_3),
    .io_mem_input_bits_4(router_io_mem_input_bits_4),
    .io_mem_input_bits_5(router_io_mem_input_bits_5),
    .io_mem_input_bits_6(router_io_mem_input_bits_6),
    .io_mem_input_bits_7(router_io_mem_input_bits_7),
    .io_mem_input_bits_8(router_io_mem_input_bits_8),
    .io_mem_input_bits_9(router_io_mem_input_bits_9),
    .io_mem_input_bits_10(router_io_mem_input_bits_10),
    .io_mem_input_bits_11(router_io_mem_input_bits_11),
    .io_mem_input_bits_12(router_io_mem_input_bits_12),
    .io_mem_input_bits_13(router_io_mem_input_bits_13),
    .io_mem_input_bits_14(router_io_mem_input_bits_14),
    .io_mem_input_bits_15(router_io_mem_input_bits_15),
    .io_mem_input_bits_16(router_io_mem_input_bits_16),
    .io_mem_input_bits_17(router_io_mem_input_bits_17),
    .io_mem_input_bits_18(router_io_mem_input_bits_18),
    .io_mem_input_bits_19(router_io_mem_input_bits_19),
    .io_mem_input_bits_20(router_io_mem_input_bits_20),
    .io_mem_input_bits_21(router_io_mem_input_bits_21),
    .io_mem_input_bits_22(router_io_mem_input_bits_22),
    .io_mem_input_bits_23(router_io_mem_input_bits_23),
    .io_mem_input_bits_24(router_io_mem_input_bits_24),
    .io_mem_input_bits_25(router_io_mem_input_bits_25),
    .io_mem_input_bits_26(router_io_mem_input_bits_26),
    .io_mem_input_bits_27(router_io_mem_input_bits_27),
    .io_mem_input_bits_28(router_io_mem_input_bits_28),
    .io_mem_input_bits_29(router_io_mem_input_bits_29),
    .io_mem_input_bits_30(router_io_mem_input_bits_30),
    .io_mem_input_bits_31(router_io_mem_input_bits_31),
    .io_array_input_ready(router_io_array_input_ready),
    .io_array_input_valid(router_io_array_input_valid),
    .io_array_input_bits_0(router_io_array_input_bits_0),
    .io_array_input_bits_1(router_io_array_input_bits_1),
    .io_array_input_bits_2(router_io_array_input_bits_2),
    .io_array_input_bits_3(router_io_array_input_bits_3),
    .io_array_input_bits_4(router_io_array_input_bits_4),
    .io_array_input_bits_5(router_io_array_input_bits_5),
    .io_array_input_bits_6(router_io_array_input_bits_6),
    .io_array_input_bits_7(router_io_array_input_bits_7),
    .io_array_input_bits_8(router_io_array_input_bits_8),
    .io_array_input_bits_9(router_io_array_input_bits_9),
    .io_array_input_bits_10(router_io_array_input_bits_10),
    .io_array_input_bits_11(router_io_array_input_bits_11),
    .io_array_input_bits_12(router_io_array_input_bits_12),
    .io_array_input_bits_13(router_io_array_input_bits_13),
    .io_array_input_bits_14(router_io_array_input_bits_14),
    .io_array_input_bits_15(router_io_array_input_bits_15),
    .io_array_input_bits_16(router_io_array_input_bits_16),
    .io_array_input_bits_17(router_io_array_input_bits_17),
    .io_array_input_bits_18(router_io_array_input_bits_18),
    .io_array_input_bits_19(router_io_array_input_bits_19),
    .io_array_input_bits_20(router_io_array_input_bits_20),
    .io_array_input_bits_21(router_io_array_input_bits_21),
    .io_array_input_bits_22(router_io_array_input_bits_22),
    .io_array_input_bits_23(router_io_array_input_bits_23),
    .io_array_input_bits_24(router_io_array_input_bits_24),
    .io_array_input_bits_25(router_io_array_input_bits_25),
    .io_array_input_bits_26(router_io_array_input_bits_26),
    .io_array_input_bits_27(router_io_array_input_bits_27),
    .io_array_input_bits_28(router_io_array_input_bits_28),
    .io_array_input_bits_29(router_io_array_input_bits_29),
    .io_array_input_bits_30(router_io_array_input_bits_30),
    .io_array_input_bits_31(router_io_array_input_bits_31),
    .io_array_output_ready(router_io_array_output_ready),
    .io_array_output_valid(router_io_array_output_valid),
    .io_array_output_bits_0(router_io_array_output_bits_0),
    .io_array_output_bits_1(router_io_array_output_bits_1),
    .io_array_output_bits_2(router_io_array_output_bits_2),
    .io_array_output_bits_3(router_io_array_output_bits_3),
    .io_array_output_bits_4(router_io_array_output_bits_4),
    .io_array_output_bits_5(router_io_array_output_bits_5),
    .io_array_output_bits_6(router_io_array_output_bits_6),
    .io_array_output_bits_7(router_io_array_output_bits_7),
    .io_array_output_bits_8(router_io_array_output_bits_8),
    .io_array_output_bits_9(router_io_array_output_bits_9),
    .io_array_output_bits_10(router_io_array_output_bits_10),
    .io_array_output_bits_11(router_io_array_output_bits_11),
    .io_array_output_bits_12(router_io_array_output_bits_12),
    .io_array_output_bits_13(router_io_array_output_bits_13),
    .io_array_output_bits_14(router_io_array_output_bits_14),
    .io_array_output_bits_15(router_io_array_output_bits_15),
    .io_array_output_bits_16(router_io_array_output_bits_16),
    .io_array_output_bits_17(router_io_array_output_bits_17),
    .io_array_output_bits_18(router_io_array_output_bits_18),
    .io_array_output_bits_19(router_io_array_output_bits_19),
    .io_array_output_bits_20(router_io_array_output_bits_20),
    .io_array_output_bits_21(router_io_array_output_bits_21),
    .io_array_output_bits_22(router_io_array_output_bits_22),
    .io_array_output_bits_23(router_io_array_output_bits_23),
    .io_array_output_bits_24(router_io_array_output_bits_24),
    .io_array_output_bits_25(router_io_array_output_bits_25),
    .io_array_output_bits_26(router_io_array_output_bits_26),
    .io_array_output_bits_27(router_io_array_output_bits_27),
    .io_array_output_bits_28(router_io_array_output_bits_28),
    .io_array_output_bits_29(router_io_array_output_bits_29),
    .io_array_output_bits_30(router_io_array_output_bits_30),
    .io_array_output_bits_31(router_io_array_output_bits_31),
    .io_array_weightInput_ready(router_io_array_weightInput_ready),
    .io_array_weightInput_valid(router_io_array_weightInput_valid),
    .io_array_weightInput_bits_0(router_io_array_weightInput_bits_0),
    .io_array_weightInput_bits_1(router_io_array_weightInput_bits_1),
    .io_array_weightInput_bits_2(router_io_array_weightInput_bits_2),
    .io_array_weightInput_bits_3(router_io_array_weightInput_bits_3),
    .io_array_weightInput_bits_4(router_io_array_weightInput_bits_4),
    .io_array_weightInput_bits_5(router_io_array_weightInput_bits_5),
    .io_array_weightInput_bits_6(router_io_array_weightInput_bits_6),
    .io_array_weightInput_bits_7(router_io_array_weightInput_bits_7),
    .io_array_weightInput_bits_8(router_io_array_weightInput_bits_8),
    .io_array_weightInput_bits_9(router_io_array_weightInput_bits_9),
    .io_array_weightInput_bits_10(router_io_array_weightInput_bits_10),
    .io_array_weightInput_bits_11(router_io_array_weightInput_bits_11),
    .io_array_weightInput_bits_12(router_io_array_weightInput_bits_12),
    .io_array_weightInput_bits_13(router_io_array_weightInput_bits_13),
    .io_array_weightInput_bits_14(router_io_array_weightInput_bits_14),
    .io_array_weightInput_bits_15(router_io_array_weightInput_bits_15),
    .io_array_weightInput_bits_16(router_io_array_weightInput_bits_16),
    .io_array_weightInput_bits_17(router_io_array_weightInput_bits_17),
    .io_array_weightInput_bits_18(router_io_array_weightInput_bits_18),
    .io_array_weightInput_bits_19(router_io_array_weightInput_bits_19),
    .io_array_weightInput_bits_20(router_io_array_weightInput_bits_20),
    .io_array_weightInput_bits_21(router_io_array_weightInput_bits_21),
    .io_array_weightInput_bits_22(router_io_array_weightInput_bits_22),
    .io_array_weightInput_bits_23(router_io_array_weightInput_bits_23),
    .io_array_weightInput_bits_24(router_io_array_weightInput_bits_24),
    .io_array_weightInput_bits_25(router_io_array_weightInput_bits_25),
    .io_array_weightInput_bits_26(router_io_array_weightInput_bits_26),
    .io_array_weightInput_bits_27(router_io_array_weightInput_bits_27),
    .io_array_weightInput_bits_28(router_io_array_weightInput_bits_28),
    .io_array_weightInput_bits_29(router_io_array_weightInput_bits_29),
    .io_array_weightInput_bits_30(router_io_array_weightInput_bits_30),
    .io_array_weightInput_bits_31(router_io_array_weightInput_bits_31),
    .io_acc_output_ready(router_io_acc_output_ready),
    .io_acc_output_valid(router_io_acc_output_valid),
    .io_acc_output_bits_0(router_io_acc_output_bits_0),
    .io_acc_output_bits_1(router_io_acc_output_bits_1),
    .io_acc_output_bits_2(router_io_acc_output_bits_2),
    .io_acc_output_bits_3(router_io_acc_output_bits_3),
    .io_acc_output_bits_4(router_io_acc_output_bits_4),
    .io_acc_output_bits_5(router_io_acc_output_bits_5),
    .io_acc_output_bits_6(router_io_acc_output_bits_6),
    .io_acc_output_bits_7(router_io_acc_output_bits_7),
    .io_acc_output_bits_8(router_io_acc_output_bits_8),
    .io_acc_output_bits_9(router_io_acc_output_bits_9),
    .io_acc_output_bits_10(router_io_acc_output_bits_10),
    .io_acc_output_bits_11(router_io_acc_output_bits_11),
    .io_acc_output_bits_12(router_io_acc_output_bits_12),
    .io_acc_output_bits_13(router_io_acc_output_bits_13),
    .io_acc_output_bits_14(router_io_acc_output_bits_14),
    .io_acc_output_bits_15(router_io_acc_output_bits_15),
    .io_acc_output_bits_16(router_io_acc_output_bits_16),
    .io_acc_output_bits_17(router_io_acc_output_bits_17),
    .io_acc_output_bits_18(router_io_acc_output_bits_18),
    .io_acc_output_bits_19(router_io_acc_output_bits_19),
    .io_acc_output_bits_20(router_io_acc_output_bits_20),
    .io_acc_output_bits_21(router_io_acc_output_bits_21),
    .io_acc_output_bits_22(router_io_acc_output_bits_22),
    .io_acc_output_bits_23(router_io_acc_output_bits_23),
    .io_acc_output_bits_24(router_io_acc_output_bits_24),
    .io_acc_output_bits_25(router_io_acc_output_bits_25),
    .io_acc_output_bits_26(router_io_acc_output_bits_26),
    .io_acc_output_bits_27(router_io_acc_output_bits_27),
    .io_acc_output_bits_28(router_io_acc_output_bits_28),
    .io_acc_output_bits_29(router_io_acc_output_bits_29),
    .io_acc_output_bits_30(router_io_acc_output_bits_30),
    .io_acc_output_bits_31(router_io_acc_output_bits_31),
    .io_acc_input_ready(router_io_acc_input_ready),
    .io_acc_input_valid(router_io_acc_input_valid),
    .io_acc_input_bits_0(router_io_acc_input_bits_0),
    .io_acc_input_bits_1(router_io_acc_input_bits_1),
    .io_acc_input_bits_2(router_io_acc_input_bits_2),
    .io_acc_input_bits_3(router_io_acc_input_bits_3),
    .io_acc_input_bits_4(router_io_acc_input_bits_4),
    .io_acc_input_bits_5(router_io_acc_input_bits_5),
    .io_acc_input_bits_6(router_io_acc_input_bits_6),
    .io_acc_input_bits_7(router_io_acc_input_bits_7),
    .io_acc_input_bits_8(router_io_acc_input_bits_8),
    .io_acc_input_bits_9(router_io_acc_input_bits_9),
    .io_acc_input_bits_10(router_io_acc_input_bits_10),
    .io_acc_input_bits_11(router_io_acc_input_bits_11),
    .io_acc_input_bits_12(router_io_acc_input_bits_12),
    .io_acc_input_bits_13(router_io_acc_input_bits_13),
    .io_acc_input_bits_14(router_io_acc_input_bits_14),
    .io_acc_input_bits_15(router_io_acc_input_bits_15),
    .io_acc_input_bits_16(router_io_acc_input_bits_16),
    .io_acc_input_bits_17(router_io_acc_input_bits_17),
    .io_acc_input_bits_18(router_io_acc_input_bits_18),
    .io_acc_input_bits_19(router_io_acc_input_bits_19),
    .io_acc_input_bits_20(router_io_acc_input_bits_20),
    .io_acc_input_bits_21(router_io_acc_input_bits_21),
    .io_acc_input_bits_22(router_io_acc_input_bits_22),
    .io_acc_input_bits_23(router_io_acc_input_bits_23),
    .io_acc_input_bits_24(router_io_acc_input_bits_24),
    .io_acc_input_bits_25(router_io_acc_input_bits_25),
    .io_acc_input_bits_26(router_io_acc_input_bits_26),
    .io_acc_input_bits_27(router_io_acc_input_bits_27),
    .io_acc_input_bits_28(router_io_acc_input_bits_28),
    .io_acc_input_bits_29(router_io_acc_input_bits_29),
    .io_acc_input_bits_30(router_io_acc_input_bits_30),
    .io_acc_input_bits_31(router_io_acc_input_bits_31),
    .io_timeout(router_io_timeout),
    .io_tracepoint(router_io_tracepoint),
    .io_programCounter(router_io_programCounter)
  );
  HostRouter hostRouter ( // @[TCU.scala 87:26]
    .io_control_ready(hostRouter_io_control_ready),
    .io_control_valid(hostRouter_io_control_valid),
    .io_control_bits_kind(hostRouter_io_control_bits_kind),
    .io_dram0_dataIn_ready(hostRouter_io_dram0_dataIn_ready),
    .io_dram0_dataIn_valid(hostRouter_io_dram0_dataIn_valid),
    .io_dram0_dataIn_bits_0(hostRouter_io_dram0_dataIn_bits_0),
    .io_dram0_dataIn_bits_1(hostRouter_io_dram0_dataIn_bits_1),
    .io_dram0_dataIn_bits_2(hostRouter_io_dram0_dataIn_bits_2),
    .io_dram0_dataIn_bits_3(hostRouter_io_dram0_dataIn_bits_3),
    .io_dram0_dataIn_bits_4(hostRouter_io_dram0_dataIn_bits_4),
    .io_dram0_dataIn_bits_5(hostRouter_io_dram0_dataIn_bits_5),
    .io_dram0_dataIn_bits_6(hostRouter_io_dram0_dataIn_bits_6),
    .io_dram0_dataIn_bits_7(hostRouter_io_dram0_dataIn_bits_7),
    .io_dram0_dataIn_bits_8(hostRouter_io_dram0_dataIn_bits_8),
    .io_dram0_dataIn_bits_9(hostRouter_io_dram0_dataIn_bits_9),
    .io_dram0_dataIn_bits_10(hostRouter_io_dram0_dataIn_bits_10),
    .io_dram0_dataIn_bits_11(hostRouter_io_dram0_dataIn_bits_11),
    .io_dram0_dataIn_bits_12(hostRouter_io_dram0_dataIn_bits_12),
    .io_dram0_dataIn_bits_13(hostRouter_io_dram0_dataIn_bits_13),
    .io_dram0_dataIn_bits_14(hostRouter_io_dram0_dataIn_bits_14),
    .io_dram0_dataIn_bits_15(hostRouter_io_dram0_dataIn_bits_15),
    .io_dram0_dataIn_bits_16(hostRouter_io_dram0_dataIn_bits_16),
    .io_dram0_dataIn_bits_17(hostRouter_io_dram0_dataIn_bits_17),
    .io_dram0_dataIn_bits_18(hostRouter_io_dram0_dataIn_bits_18),
    .io_dram0_dataIn_bits_19(hostRouter_io_dram0_dataIn_bits_19),
    .io_dram0_dataIn_bits_20(hostRouter_io_dram0_dataIn_bits_20),
    .io_dram0_dataIn_bits_21(hostRouter_io_dram0_dataIn_bits_21),
    .io_dram0_dataIn_bits_22(hostRouter_io_dram0_dataIn_bits_22),
    .io_dram0_dataIn_bits_23(hostRouter_io_dram0_dataIn_bits_23),
    .io_dram0_dataIn_bits_24(hostRouter_io_dram0_dataIn_bits_24),
    .io_dram0_dataIn_bits_25(hostRouter_io_dram0_dataIn_bits_25),
    .io_dram0_dataIn_bits_26(hostRouter_io_dram0_dataIn_bits_26),
    .io_dram0_dataIn_bits_27(hostRouter_io_dram0_dataIn_bits_27),
    .io_dram0_dataIn_bits_28(hostRouter_io_dram0_dataIn_bits_28),
    .io_dram0_dataIn_bits_29(hostRouter_io_dram0_dataIn_bits_29),
    .io_dram0_dataIn_bits_30(hostRouter_io_dram0_dataIn_bits_30),
    .io_dram0_dataIn_bits_31(hostRouter_io_dram0_dataIn_bits_31),
    .io_dram0_dataOut_ready(hostRouter_io_dram0_dataOut_ready),
    .io_dram0_dataOut_valid(hostRouter_io_dram0_dataOut_valid),
    .io_dram0_dataOut_bits_0(hostRouter_io_dram0_dataOut_bits_0),
    .io_dram0_dataOut_bits_1(hostRouter_io_dram0_dataOut_bits_1),
    .io_dram0_dataOut_bits_2(hostRouter_io_dram0_dataOut_bits_2),
    .io_dram0_dataOut_bits_3(hostRouter_io_dram0_dataOut_bits_3),
    .io_dram0_dataOut_bits_4(hostRouter_io_dram0_dataOut_bits_4),
    .io_dram0_dataOut_bits_5(hostRouter_io_dram0_dataOut_bits_5),
    .io_dram0_dataOut_bits_6(hostRouter_io_dram0_dataOut_bits_6),
    .io_dram0_dataOut_bits_7(hostRouter_io_dram0_dataOut_bits_7),
    .io_dram0_dataOut_bits_8(hostRouter_io_dram0_dataOut_bits_8),
    .io_dram0_dataOut_bits_9(hostRouter_io_dram0_dataOut_bits_9),
    .io_dram0_dataOut_bits_10(hostRouter_io_dram0_dataOut_bits_10),
    .io_dram0_dataOut_bits_11(hostRouter_io_dram0_dataOut_bits_11),
    .io_dram0_dataOut_bits_12(hostRouter_io_dram0_dataOut_bits_12),
    .io_dram0_dataOut_bits_13(hostRouter_io_dram0_dataOut_bits_13),
    .io_dram0_dataOut_bits_14(hostRouter_io_dram0_dataOut_bits_14),
    .io_dram0_dataOut_bits_15(hostRouter_io_dram0_dataOut_bits_15),
    .io_dram0_dataOut_bits_16(hostRouter_io_dram0_dataOut_bits_16),
    .io_dram0_dataOut_bits_17(hostRouter_io_dram0_dataOut_bits_17),
    .io_dram0_dataOut_bits_18(hostRouter_io_dram0_dataOut_bits_18),
    .io_dram0_dataOut_bits_19(hostRouter_io_dram0_dataOut_bits_19),
    .io_dram0_dataOut_bits_20(hostRouter_io_dram0_dataOut_bits_20),
    .io_dram0_dataOut_bits_21(hostRouter_io_dram0_dataOut_bits_21),
    .io_dram0_dataOut_bits_22(hostRouter_io_dram0_dataOut_bits_22),
    .io_dram0_dataOut_bits_23(hostRouter_io_dram0_dataOut_bits_23),
    .io_dram0_dataOut_bits_24(hostRouter_io_dram0_dataOut_bits_24),
    .io_dram0_dataOut_bits_25(hostRouter_io_dram0_dataOut_bits_25),
    .io_dram0_dataOut_bits_26(hostRouter_io_dram0_dataOut_bits_26),
    .io_dram0_dataOut_bits_27(hostRouter_io_dram0_dataOut_bits_27),
    .io_dram0_dataOut_bits_28(hostRouter_io_dram0_dataOut_bits_28),
    .io_dram0_dataOut_bits_29(hostRouter_io_dram0_dataOut_bits_29),
    .io_dram0_dataOut_bits_30(hostRouter_io_dram0_dataOut_bits_30),
    .io_dram0_dataOut_bits_31(hostRouter_io_dram0_dataOut_bits_31),
    .io_dram1_dataIn_ready(hostRouter_io_dram1_dataIn_ready),
    .io_dram1_dataIn_valid(hostRouter_io_dram1_dataIn_valid),
    .io_dram1_dataIn_bits_0(hostRouter_io_dram1_dataIn_bits_0),
    .io_dram1_dataIn_bits_1(hostRouter_io_dram1_dataIn_bits_1),
    .io_dram1_dataIn_bits_2(hostRouter_io_dram1_dataIn_bits_2),
    .io_dram1_dataIn_bits_3(hostRouter_io_dram1_dataIn_bits_3),
    .io_dram1_dataIn_bits_4(hostRouter_io_dram1_dataIn_bits_4),
    .io_dram1_dataIn_bits_5(hostRouter_io_dram1_dataIn_bits_5),
    .io_dram1_dataIn_bits_6(hostRouter_io_dram1_dataIn_bits_6),
    .io_dram1_dataIn_bits_7(hostRouter_io_dram1_dataIn_bits_7),
    .io_dram1_dataIn_bits_8(hostRouter_io_dram1_dataIn_bits_8),
    .io_dram1_dataIn_bits_9(hostRouter_io_dram1_dataIn_bits_9),
    .io_dram1_dataIn_bits_10(hostRouter_io_dram1_dataIn_bits_10),
    .io_dram1_dataIn_bits_11(hostRouter_io_dram1_dataIn_bits_11),
    .io_dram1_dataIn_bits_12(hostRouter_io_dram1_dataIn_bits_12),
    .io_dram1_dataIn_bits_13(hostRouter_io_dram1_dataIn_bits_13),
    .io_dram1_dataIn_bits_14(hostRouter_io_dram1_dataIn_bits_14),
    .io_dram1_dataIn_bits_15(hostRouter_io_dram1_dataIn_bits_15),
    .io_dram1_dataIn_bits_16(hostRouter_io_dram1_dataIn_bits_16),
    .io_dram1_dataIn_bits_17(hostRouter_io_dram1_dataIn_bits_17),
    .io_dram1_dataIn_bits_18(hostRouter_io_dram1_dataIn_bits_18),
    .io_dram1_dataIn_bits_19(hostRouter_io_dram1_dataIn_bits_19),
    .io_dram1_dataIn_bits_20(hostRouter_io_dram1_dataIn_bits_20),
    .io_dram1_dataIn_bits_21(hostRouter_io_dram1_dataIn_bits_21),
    .io_dram1_dataIn_bits_22(hostRouter_io_dram1_dataIn_bits_22),
    .io_dram1_dataIn_bits_23(hostRouter_io_dram1_dataIn_bits_23),
    .io_dram1_dataIn_bits_24(hostRouter_io_dram1_dataIn_bits_24),
    .io_dram1_dataIn_bits_25(hostRouter_io_dram1_dataIn_bits_25),
    .io_dram1_dataIn_bits_26(hostRouter_io_dram1_dataIn_bits_26),
    .io_dram1_dataIn_bits_27(hostRouter_io_dram1_dataIn_bits_27),
    .io_dram1_dataIn_bits_28(hostRouter_io_dram1_dataIn_bits_28),
    .io_dram1_dataIn_bits_29(hostRouter_io_dram1_dataIn_bits_29),
    .io_dram1_dataIn_bits_30(hostRouter_io_dram1_dataIn_bits_30),
    .io_dram1_dataIn_bits_31(hostRouter_io_dram1_dataIn_bits_31),
    .io_dram1_dataOut_ready(hostRouter_io_dram1_dataOut_ready),
    .io_dram1_dataOut_valid(hostRouter_io_dram1_dataOut_valid),
    .io_dram1_dataOut_bits_0(hostRouter_io_dram1_dataOut_bits_0),
    .io_dram1_dataOut_bits_1(hostRouter_io_dram1_dataOut_bits_1),
    .io_dram1_dataOut_bits_2(hostRouter_io_dram1_dataOut_bits_2),
    .io_dram1_dataOut_bits_3(hostRouter_io_dram1_dataOut_bits_3),
    .io_dram1_dataOut_bits_4(hostRouter_io_dram1_dataOut_bits_4),
    .io_dram1_dataOut_bits_5(hostRouter_io_dram1_dataOut_bits_5),
    .io_dram1_dataOut_bits_6(hostRouter_io_dram1_dataOut_bits_6),
    .io_dram1_dataOut_bits_7(hostRouter_io_dram1_dataOut_bits_7),
    .io_dram1_dataOut_bits_8(hostRouter_io_dram1_dataOut_bits_8),
    .io_dram1_dataOut_bits_9(hostRouter_io_dram1_dataOut_bits_9),
    .io_dram1_dataOut_bits_10(hostRouter_io_dram1_dataOut_bits_10),
    .io_dram1_dataOut_bits_11(hostRouter_io_dram1_dataOut_bits_11),
    .io_dram1_dataOut_bits_12(hostRouter_io_dram1_dataOut_bits_12),
    .io_dram1_dataOut_bits_13(hostRouter_io_dram1_dataOut_bits_13),
    .io_dram1_dataOut_bits_14(hostRouter_io_dram1_dataOut_bits_14),
    .io_dram1_dataOut_bits_15(hostRouter_io_dram1_dataOut_bits_15),
    .io_dram1_dataOut_bits_16(hostRouter_io_dram1_dataOut_bits_16),
    .io_dram1_dataOut_bits_17(hostRouter_io_dram1_dataOut_bits_17),
    .io_dram1_dataOut_bits_18(hostRouter_io_dram1_dataOut_bits_18),
    .io_dram1_dataOut_bits_19(hostRouter_io_dram1_dataOut_bits_19),
    .io_dram1_dataOut_bits_20(hostRouter_io_dram1_dataOut_bits_20),
    .io_dram1_dataOut_bits_21(hostRouter_io_dram1_dataOut_bits_21),
    .io_dram1_dataOut_bits_22(hostRouter_io_dram1_dataOut_bits_22),
    .io_dram1_dataOut_bits_23(hostRouter_io_dram1_dataOut_bits_23),
    .io_dram1_dataOut_bits_24(hostRouter_io_dram1_dataOut_bits_24),
    .io_dram1_dataOut_bits_25(hostRouter_io_dram1_dataOut_bits_25),
    .io_dram1_dataOut_bits_26(hostRouter_io_dram1_dataOut_bits_26),
    .io_dram1_dataOut_bits_27(hostRouter_io_dram1_dataOut_bits_27),
    .io_dram1_dataOut_bits_28(hostRouter_io_dram1_dataOut_bits_28),
    .io_dram1_dataOut_bits_29(hostRouter_io_dram1_dataOut_bits_29),
    .io_dram1_dataOut_bits_30(hostRouter_io_dram1_dataOut_bits_30),
    .io_dram1_dataOut_bits_31(hostRouter_io_dram1_dataOut_bits_31),
    .io_mem_output_ready(hostRouter_io_mem_output_ready),
    .io_mem_output_valid(hostRouter_io_mem_output_valid),
    .io_mem_output_bits_0(hostRouter_io_mem_output_bits_0),
    .io_mem_output_bits_1(hostRouter_io_mem_output_bits_1),
    .io_mem_output_bits_2(hostRouter_io_mem_output_bits_2),
    .io_mem_output_bits_3(hostRouter_io_mem_output_bits_3),
    .io_mem_output_bits_4(hostRouter_io_mem_output_bits_4),
    .io_mem_output_bits_5(hostRouter_io_mem_output_bits_5),
    .io_mem_output_bits_6(hostRouter_io_mem_output_bits_6),
    .io_mem_output_bits_7(hostRouter_io_mem_output_bits_7),
    .io_mem_output_bits_8(hostRouter_io_mem_output_bits_8),
    .io_mem_output_bits_9(hostRouter_io_mem_output_bits_9),
    .io_mem_output_bits_10(hostRouter_io_mem_output_bits_10),
    .io_mem_output_bits_11(hostRouter_io_mem_output_bits_11),
    .io_mem_output_bits_12(hostRouter_io_mem_output_bits_12),
    .io_mem_output_bits_13(hostRouter_io_mem_output_bits_13),
    .io_mem_output_bits_14(hostRouter_io_mem_output_bits_14),
    .io_mem_output_bits_15(hostRouter_io_mem_output_bits_15),
    .io_mem_output_bits_16(hostRouter_io_mem_output_bits_16),
    .io_mem_output_bits_17(hostRouter_io_mem_output_bits_17),
    .io_mem_output_bits_18(hostRouter_io_mem_output_bits_18),
    .io_mem_output_bits_19(hostRouter_io_mem_output_bits_19),
    .io_mem_output_bits_20(hostRouter_io_mem_output_bits_20),
    .io_mem_output_bits_21(hostRouter_io_mem_output_bits_21),
    .io_mem_output_bits_22(hostRouter_io_mem_output_bits_22),
    .io_mem_output_bits_23(hostRouter_io_mem_output_bits_23),
    .io_mem_output_bits_24(hostRouter_io_mem_output_bits_24),
    .io_mem_output_bits_25(hostRouter_io_mem_output_bits_25),
    .io_mem_output_bits_26(hostRouter_io_mem_output_bits_26),
    .io_mem_output_bits_27(hostRouter_io_mem_output_bits_27),
    .io_mem_output_bits_28(hostRouter_io_mem_output_bits_28),
    .io_mem_output_bits_29(hostRouter_io_mem_output_bits_29),
    .io_mem_output_bits_30(hostRouter_io_mem_output_bits_30),
    .io_mem_output_bits_31(hostRouter_io_mem_output_bits_31),
    .io_mem_input_ready(hostRouter_io_mem_input_ready),
    .io_mem_input_valid(hostRouter_io_mem_input_valid),
    .io_mem_input_bits_0(hostRouter_io_mem_input_bits_0),
    .io_mem_input_bits_1(hostRouter_io_mem_input_bits_1),
    .io_mem_input_bits_2(hostRouter_io_mem_input_bits_2),
    .io_mem_input_bits_3(hostRouter_io_mem_input_bits_3),
    .io_mem_input_bits_4(hostRouter_io_mem_input_bits_4),
    .io_mem_input_bits_5(hostRouter_io_mem_input_bits_5),
    .io_mem_input_bits_6(hostRouter_io_mem_input_bits_6),
    .io_mem_input_bits_7(hostRouter_io_mem_input_bits_7),
    .io_mem_input_bits_8(hostRouter_io_mem_input_bits_8),
    .io_mem_input_bits_9(hostRouter_io_mem_input_bits_9),
    .io_mem_input_bits_10(hostRouter_io_mem_input_bits_10),
    .io_mem_input_bits_11(hostRouter_io_mem_input_bits_11),
    .io_mem_input_bits_12(hostRouter_io_mem_input_bits_12),
    .io_mem_input_bits_13(hostRouter_io_mem_input_bits_13),
    .io_mem_input_bits_14(hostRouter_io_mem_input_bits_14),
    .io_mem_input_bits_15(hostRouter_io_mem_input_bits_15),
    .io_mem_input_bits_16(hostRouter_io_mem_input_bits_16),
    .io_mem_input_bits_17(hostRouter_io_mem_input_bits_17),
    .io_mem_input_bits_18(hostRouter_io_mem_input_bits_18),
    .io_mem_input_bits_19(hostRouter_io_mem_input_bits_19),
    .io_mem_input_bits_20(hostRouter_io_mem_input_bits_20),
    .io_mem_input_bits_21(hostRouter_io_mem_input_bits_21),
    .io_mem_input_bits_22(hostRouter_io_mem_input_bits_22),
    .io_mem_input_bits_23(hostRouter_io_mem_input_bits_23),
    .io_mem_input_bits_24(hostRouter_io_mem_input_bits_24),
    .io_mem_input_bits_25(hostRouter_io_mem_input_bits_25),
    .io_mem_input_bits_26(hostRouter_io_mem_input_bits_26),
    .io_mem_input_bits_27(hostRouter_io_mem_input_bits_27),
    .io_mem_input_bits_28(hostRouter_io_mem_input_bits_28),
    .io_mem_input_bits_29(hostRouter_io_mem_input_bits_29),
    .io_mem_input_bits_30(hostRouter_io_mem_input_bits_30),
    .io_mem_input_bits_31(hostRouter_io_mem_input_bits_31)
  );
  Queue_28 acc_io_control_q ( // @[TCU.scala 110:39]
    .clock(acc_io_control_q_clock),
    .reset(acc_io_control_q_reset),
    .io_enq_ready(acc_io_control_q_io_enq_ready),
    .io_enq_valid(acc_io_control_q_io_enq_valid),
    .io_enq_bits_instruction_op(acc_io_control_q_io_enq_bits_instruction_op),
    .io_enq_bits_instruction_sourceLeft(acc_io_control_q_io_enq_bits_instruction_sourceLeft),
    .io_enq_bits_instruction_sourceRight(acc_io_control_q_io_enq_bits_instruction_sourceRight),
    .io_enq_bits_instruction_dest(acc_io_control_q_io_enq_bits_instruction_dest),
    .io_enq_bits_readAddress(acc_io_control_q_io_enq_bits_readAddress),
    .io_enq_bits_writeAddress(acc_io_control_q_io_enq_bits_writeAddress),
    .io_enq_bits_accumulate(acc_io_control_q_io_enq_bits_accumulate),
    .io_enq_bits_write(acc_io_control_q_io_enq_bits_write),
    .io_enq_bits_read(acc_io_control_q_io_enq_bits_read),
    .io_deq_ready(acc_io_control_q_io_deq_ready),
    .io_deq_valid(acc_io_control_q_io_deq_valid),
    .io_deq_bits_instruction_op(acc_io_control_q_io_deq_bits_instruction_op),
    .io_deq_bits_instruction_sourceLeft(acc_io_control_q_io_deq_bits_instruction_sourceLeft),
    .io_deq_bits_instruction_sourceRight(acc_io_control_q_io_deq_bits_instruction_sourceRight),
    .io_deq_bits_instruction_dest(acc_io_control_q_io_deq_bits_instruction_dest),
    .io_deq_bits_readAddress(acc_io_control_q_io_deq_bits_readAddress),
    .io_deq_bits_writeAddress(acc_io_control_q_io_deq_bits_writeAddress),
    .io_deq_bits_accumulate(acc_io_control_q_io_deq_bits_accumulate),
    .io_deq_bits_write(acc_io_control_q_io_deq_bits_write),
    .io_deq_bits_read(acc_io_control_q_io_deq_bits_read)
  );
  Queue_29 array_io_control_q ( // @[TCU.scala 117:41]
    .clock(array_io_control_q_clock),
    .reset(array_io_control_q_reset),
    .io_enq_ready(array_io_control_q_io_enq_ready),
    .io_enq_valid(array_io_control_q_io_enq_valid),
    .io_enq_bits_load(array_io_control_q_io_enq_bits_load),
    .io_enq_bits_zeroes(array_io_control_q_io_enq_bits_zeroes),
    .io_deq_ready(array_io_control_q_io_deq_ready),
    .io_deq_valid(array_io_control_q_io_deq_valid),
    .io_deq_bits_load(array_io_control_q_io_deq_bits_load),
    .io_deq_bits_zeroes(array_io_control_q_io_deq_bits_zeroes)
  );
  assign io_instruction_ready = decoder_io_instruction_ready; // @[TCU.scala 97:26]
  assign io_dram0_control_valid = decoder_io_dram0_valid; // @[TCU.scala 99:20]
  assign io_dram0_control_bits_write = decoder_io_dram0_bits_write; // @[TCU.scala 99:20]
  assign io_dram0_control_bits_address = decoder_io_dram0_bits_address; // @[TCU.scala 99:20]
  assign io_dram0_control_bits_size = decoder_io_dram0_bits_size; // @[TCU.scala 99:20]
  assign io_dram0_dataIn_ready = hostRouter_io_dram0_dataIn_ready; // @[TCU.scala 155:30]
  assign io_dram0_dataOut_valid = hostRouter_io_dram0_dataOut_valid; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_0 = hostRouter_io_dram0_dataOut_bits_0; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_1 = hostRouter_io_dram0_dataOut_bits_1; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_2 = hostRouter_io_dram0_dataOut_bits_2; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_3 = hostRouter_io_dram0_dataOut_bits_3; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_4 = hostRouter_io_dram0_dataOut_bits_4; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_5 = hostRouter_io_dram0_dataOut_bits_5; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_6 = hostRouter_io_dram0_dataOut_bits_6; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_7 = hostRouter_io_dram0_dataOut_bits_7; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_8 = hostRouter_io_dram0_dataOut_bits_8; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_9 = hostRouter_io_dram0_dataOut_bits_9; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_10 = hostRouter_io_dram0_dataOut_bits_10; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_11 = hostRouter_io_dram0_dataOut_bits_11; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_12 = hostRouter_io_dram0_dataOut_bits_12; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_13 = hostRouter_io_dram0_dataOut_bits_13; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_14 = hostRouter_io_dram0_dataOut_bits_14; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_15 = hostRouter_io_dram0_dataOut_bits_15; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_16 = hostRouter_io_dram0_dataOut_bits_16; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_17 = hostRouter_io_dram0_dataOut_bits_17; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_18 = hostRouter_io_dram0_dataOut_bits_18; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_19 = hostRouter_io_dram0_dataOut_bits_19; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_20 = hostRouter_io_dram0_dataOut_bits_20; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_21 = hostRouter_io_dram0_dataOut_bits_21; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_22 = hostRouter_io_dram0_dataOut_bits_22; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_23 = hostRouter_io_dram0_dataOut_bits_23; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_24 = hostRouter_io_dram0_dataOut_bits_24; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_25 = hostRouter_io_dram0_dataOut_bits_25; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_26 = hostRouter_io_dram0_dataOut_bits_26; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_27 = hostRouter_io_dram0_dataOut_bits_27; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_28 = hostRouter_io_dram0_dataOut_bits_28; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_29 = hostRouter_io_dram0_dataOut_bits_29; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_30 = hostRouter_io_dram0_dataOut_bits_30; // @[TCU.scala 156:20]
  assign io_dram0_dataOut_bits_31 = hostRouter_io_dram0_dataOut_bits_31; // @[TCU.scala 156:20]
  assign io_dram1_control_valid = decoder_io_dram1_valid; // @[TCU.scala 100:20]
  assign io_dram1_control_bits_write = decoder_io_dram1_bits_write; // @[TCU.scala 100:20]
  assign io_dram1_control_bits_address = decoder_io_dram1_bits_address; // @[TCU.scala 100:20]
  assign io_dram1_control_bits_size = decoder_io_dram1_bits_size; // @[TCU.scala 100:20]
  assign io_dram1_dataIn_ready = hostRouter_io_dram1_dataIn_ready; // @[TCU.scala 158:30]
  assign io_dram1_dataOut_valid = hostRouter_io_dram1_dataOut_valid; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_0 = hostRouter_io_dram1_dataOut_bits_0; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_1 = hostRouter_io_dram1_dataOut_bits_1; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_2 = hostRouter_io_dram1_dataOut_bits_2; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_3 = hostRouter_io_dram1_dataOut_bits_3; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_4 = hostRouter_io_dram1_dataOut_bits_4; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_5 = hostRouter_io_dram1_dataOut_bits_5; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_6 = hostRouter_io_dram1_dataOut_bits_6; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_7 = hostRouter_io_dram1_dataOut_bits_7; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_8 = hostRouter_io_dram1_dataOut_bits_8; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_9 = hostRouter_io_dram1_dataOut_bits_9; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_10 = hostRouter_io_dram1_dataOut_bits_10; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_11 = hostRouter_io_dram1_dataOut_bits_11; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_12 = hostRouter_io_dram1_dataOut_bits_12; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_13 = hostRouter_io_dram1_dataOut_bits_13; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_14 = hostRouter_io_dram1_dataOut_bits_14; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_15 = hostRouter_io_dram1_dataOut_bits_15; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_16 = hostRouter_io_dram1_dataOut_bits_16; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_17 = hostRouter_io_dram1_dataOut_bits_17; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_18 = hostRouter_io_dram1_dataOut_bits_18; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_19 = hostRouter_io_dram1_dataOut_bits_19; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_20 = hostRouter_io_dram1_dataOut_bits_20; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_21 = hostRouter_io_dram1_dataOut_bits_21; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_22 = hostRouter_io_dram1_dataOut_bits_22; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_23 = hostRouter_io_dram1_dataOut_bits_23; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_24 = hostRouter_io_dram1_dataOut_bits_24; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_25 = hostRouter_io_dram1_dataOut_bits_25; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_26 = hostRouter_io_dram1_dataOut_bits_26; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_27 = hostRouter_io_dram1_dataOut_bits_27; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_28 = hostRouter_io_dram1_dataOut_bits_28; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_29 = hostRouter_io_dram1_dataOut_bits_29; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_30 = hostRouter_io_dram1_dataOut_bits_30; // @[TCU.scala 159:20]
  assign io_dram1_dataOut_bits_31 = hostRouter_io_dram1_dataOut_bits_31; // @[TCU.scala 159:20]
  assign io_config_dram0AddressOffset = decoder_io_config_dram0AddressOffset; // @[TCU.scala 101:13]
  assign io_config_dram0CacheBehaviour = decoder_io_config_dram0CacheBehaviour; // @[TCU.scala 101:13]
  assign io_config_dram1AddressOffset = decoder_io_config_dram1AddressOffset; // @[TCU.scala 101:13]
  assign io_config_dram1CacheBehaviour = decoder_io_config_dram1CacheBehaviour; // @[TCU.scala 101:13]
  assign io_timeout = decoder_io_timeout; // @[TCU.scala 102:14]
  assign io_tracepoint = decoder_io_tracepoint; // @[TCU.scala 104:17]
  assign io_programCounter = decoder_io_programCounter; // @[TCU.scala 105:21]
  assign decoder_clock = clock;
  assign decoder_reset = reset;
  assign decoder_io_instruction_valid = io_instruction_valid; // @[TCU.scala 97:26]
  assign decoder_io_instruction_bits_opcode = io_instruction_bits_opcode; // @[TCU.scala 97:26]
  assign decoder_io_instruction_bits_flags = io_instruction_bits_flags; // @[TCU.scala 97:26]
  assign decoder_io_instruction_bits_arguments = io_instruction_bits_arguments; // @[TCU.scala 97:26]
  assign decoder_io_memPortA_ready = mem_io_portA_control_ready; // @[TCU.scala 124:17]
  assign decoder_io_memPortB_ready = mem_io_portB_control_ready; // @[TCU.scala 148:17]
  assign decoder_io_dram0_ready = io_dram0_control_ready; // @[TCU.scala 99:20]
  assign decoder_io_dram1_ready = io_dram1_control_ready; // @[TCU.scala 100:20]
  assign decoder_io_dataflow_ready = router_io_control_ready; // @[TCU.scala 133:21]
  assign decoder_io_hostDataflow_ready = hostRouter_io_control_ready; // @[TCU.scala 146:25]
  assign decoder_io_acc_ready = acc_io_control_q_io_enq_ready; // @[TCU.scala 110:39]
  assign decoder_io_array_ready = array_io_control_q_io_enq_ready; // @[TCU.scala 117:41]
  assign array_clock = clock;
  assign array_reset = reset;
  assign array_io_control_valid = array_io_control_q_io_deq_valid; // @[TCU.scala 117:20]
  assign array_io_control_bits_load = array_io_control_q_io_deq_bits_load; // @[TCU.scala 117:20]
  assign array_io_control_bits_zeroes = array_io_control_q_io_deq_bits_zeroes; // @[TCU.scala 117:20]
  assign array_io_input_valid = router_io_array_input_valid; // @[TCU.scala 138:18]
  assign array_io_input_bits_0 = router_io_array_input_bits_0; // @[TCU.scala 138:18]
  assign array_io_input_bits_1 = router_io_array_input_bits_1; // @[TCU.scala 138:18]
  assign array_io_input_bits_2 = router_io_array_input_bits_2; // @[TCU.scala 138:18]
  assign array_io_input_bits_3 = router_io_array_input_bits_3; // @[TCU.scala 138:18]
  assign array_io_input_bits_4 = router_io_array_input_bits_4; // @[TCU.scala 138:18]
  assign array_io_input_bits_5 = router_io_array_input_bits_5; // @[TCU.scala 138:18]
  assign array_io_input_bits_6 = router_io_array_input_bits_6; // @[TCU.scala 138:18]
  assign array_io_input_bits_7 = router_io_array_input_bits_7; // @[TCU.scala 138:18]
  assign array_io_input_bits_8 = router_io_array_input_bits_8; // @[TCU.scala 138:18]
  assign array_io_input_bits_9 = router_io_array_input_bits_9; // @[TCU.scala 138:18]
  assign array_io_input_bits_10 = router_io_array_input_bits_10; // @[TCU.scala 138:18]
  assign array_io_input_bits_11 = router_io_array_input_bits_11; // @[TCU.scala 138:18]
  assign array_io_input_bits_12 = router_io_array_input_bits_12; // @[TCU.scala 138:18]
  assign array_io_input_bits_13 = router_io_array_input_bits_13; // @[TCU.scala 138:18]
  assign array_io_input_bits_14 = router_io_array_input_bits_14; // @[TCU.scala 138:18]
  assign array_io_input_bits_15 = router_io_array_input_bits_15; // @[TCU.scala 138:18]
  assign array_io_input_bits_16 = router_io_array_input_bits_16; // @[TCU.scala 138:18]
  assign array_io_input_bits_17 = router_io_array_input_bits_17; // @[TCU.scala 138:18]
  assign array_io_input_bits_18 = router_io_array_input_bits_18; // @[TCU.scala 138:18]
  assign array_io_input_bits_19 = router_io_array_input_bits_19; // @[TCU.scala 138:18]
  assign array_io_input_bits_20 = router_io_array_input_bits_20; // @[TCU.scala 138:18]
  assign array_io_input_bits_21 = router_io_array_input_bits_21; // @[TCU.scala 138:18]
  assign array_io_input_bits_22 = router_io_array_input_bits_22; // @[TCU.scala 138:18]
  assign array_io_input_bits_23 = router_io_array_input_bits_23; // @[TCU.scala 138:18]
  assign array_io_input_bits_24 = router_io_array_input_bits_24; // @[TCU.scala 138:18]
  assign array_io_input_bits_25 = router_io_array_input_bits_25; // @[TCU.scala 138:18]
  assign array_io_input_bits_26 = router_io_array_input_bits_26; // @[TCU.scala 138:18]
  assign array_io_input_bits_27 = router_io_array_input_bits_27; // @[TCU.scala 138:18]
  assign array_io_input_bits_28 = router_io_array_input_bits_28; // @[TCU.scala 138:18]
  assign array_io_input_bits_29 = router_io_array_input_bits_29; // @[TCU.scala 138:18]
  assign array_io_input_bits_30 = router_io_array_input_bits_30; // @[TCU.scala 138:18]
  assign array_io_input_bits_31 = router_io_array_input_bits_31; // @[TCU.scala 138:18]
  assign array_io_weight_valid = router_io_array_weightInput_valid; // @[TCU.scala 140:19]
  assign array_io_weight_bits_0 = router_io_array_weightInput_bits_0; // @[TCU.scala 140:19]
  assign array_io_weight_bits_1 = router_io_array_weightInput_bits_1; // @[TCU.scala 140:19]
  assign array_io_weight_bits_2 = router_io_array_weightInput_bits_2; // @[TCU.scala 140:19]
  assign array_io_weight_bits_3 = router_io_array_weightInput_bits_3; // @[TCU.scala 140:19]
  assign array_io_weight_bits_4 = router_io_array_weightInput_bits_4; // @[TCU.scala 140:19]
  assign array_io_weight_bits_5 = router_io_array_weightInput_bits_5; // @[TCU.scala 140:19]
  assign array_io_weight_bits_6 = router_io_array_weightInput_bits_6; // @[TCU.scala 140:19]
  assign array_io_weight_bits_7 = router_io_array_weightInput_bits_7; // @[TCU.scala 140:19]
  assign array_io_weight_bits_8 = router_io_array_weightInput_bits_8; // @[TCU.scala 140:19]
  assign array_io_weight_bits_9 = router_io_array_weightInput_bits_9; // @[TCU.scala 140:19]
  assign array_io_weight_bits_10 = router_io_array_weightInput_bits_10; // @[TCU.scala 140:19]
  assign array_io_weight_bits_11 = router_io_array_weightInput_bits_11; // @[TCU.scala 140:19]
  assign array_io_weight_bits_12 = router_io_array_weightInput_bits_12; // @[TCU.scala 140:19]
  assign array_io_weight_bits_13 = router_io_array_weightInput_bits_13; // @[TCU.scala 140:19]
  assign array_io_weight_bits_14 = router_io_array_weightInput_bits_14; // @[TCU.scala 140:19]
  assign array_io_weight_bits_15 = router_io_array_weightInput_bits_15; // @[TCU.scala 140:19]
  assign array_io_weight_bits_16 = router_io_array_weightInput_bits_16; // @[TCU.scala 140:19]
  assign array_io_weight_bits_17 = router_io_array_weightInput_bits_17; // @[TCU.scala 140:19]
  assign array_io_weight_bits_18 = router_io_array_weightInput_bits_18; // @[TCU.scala 140:19]
  assign array_io_weight_bits_19 = router_io_array_weightInput_bits_19; // @[TCU.scala 140:19]
  assign array_io_weight_bits_20 = router_io_array_weightInput_bits_20; // @[TCU.scala 140:19]
  assign array_io_weight_bits_21 = router_io_array_weightInput_bits_21; // @[TCU.scala 140:19]
  assign array_io_weight_bits_22 = router_io_array_weightInput_bits_22; // @[TCU.scala 140:19]
  assign array_io_weight_bits_23 = router_io_array_weightInput_bits_23; // @[TCU.scala 140:19]
  assign array_io_weight_bits_24 = router_io_array_weightInput_bits_24; // @[TCU.scala 140:19]
  assign array_io_weight_bits_25 = router_io_array_weightInput_bits_25; // @[TCU.scala 140:19]
  assign array_io_weight_bits_26 = router_io_array_weightInput_bits_26; // @[TCU.scala 140:19]
  assign array_io_weight_bits_27 = router_io_array_weightInput_bits_27; // @[TCU.scala 140:19]
  assign array_io_weight_bits_28 = router_io_array_weightInput_bits_28; // @[TCU.scala 140:19]
  assign array_io_weight_bits_29 = router_io_array_weightInput_bits_29; // @[TCU.scala 140:19]
  assign array_io_weight_bits_30 = router_io_array_weightInput_bits_30; // @[TCU.scala 140:19]
  assign array_io_weight_bits_31 = router_io_array_weightInput_bits_31; // @[TCU.scala 140:19]
  assign array_io_output_ready = router_io_array_output_ready; // @[TCU.scala 139:26]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_io_input_valid = router_io_acc_input_valid; // @[TCU.scala 142:16]
  assign acc_io_input_bits_0 = router_io_acc_input_bits_0; // @[TCU.scala 142:16]
  assign acc_io_input_bits_1 = router_io_acc_input_bits_1; // @[TCU.scala 142:16]
  assign acc_io_input_bits_2 = router_io_acc_input_bits_2; // @[TCU.scala 142:16]
  assign acc_io_input_bits_3 = router_io_acc_input_bits_3; // @[TCU.scala 142:16]
  assign acc_io_input_bits_4 = router_io_acc_input_bits_4; // @[TCU.scala 142:16]
  assign acc_io_input_bits_5 = router_io_acc_input_bits_5; // @[TCU.scala 142:16]
  assign acc_io_input_bits_6 = router_io_acc_input_bits_6; // @[TCU.scala 142:16]
  assign acc_io_input_bits_7 = router_io_acc_input_bits_7; // @[TCU.scala 142:16]
  assign acc_io_input_bits_8 = router_io_acc_input_bits_8; // @[TCU.scala 142:16]
  assign acc_io_input_bits_9 = router_io_acc_input_bits_9; // @[TCU.scala 142:16]
  assign acc_io_input_bits_10 = router_io_acc_input_bits_10; // @[TCU.scala 142:16]
  assign acc_io_input_bits_11 = router_io_acc_input_bits_11; // @[TCU.scala 142:16]
  assign acc_io_input_bits_12 = router_io_acc_input_bits_12; // @[TCU.scala 142:16]
  assign acc_io_input_bits_13 = router_io_acc_input_bits_13; // @[TCU.scala 142:16]
  assign acc_io_input_bits_14 = router_io_acc_input_bits_14; // @[TCU.scala 142:16]
  assign acc_io_input_bits_15 = router_io_acc_input_bits_15; // @[TCU.scala 142:16]
  assign acc_io_input_bits_16 = router_io_acc_input_bits_16; // @[TCU.scala 142:16]
  assign acc_io_input_bits_17 = router_io_acc_input_bits_17; // @[TCU.scala 142:16]
  assign acc_io_input_bits_18 = router_io_acc_input_bits_18; // @[TCU.scala 142:16]
  assign acc_io_input_bits_19 = router_io_acc_input_bits_19; // @[TCU.scala 142:16]
  assign acc_io_input_bits_20 = router_io_acc_input_bits_20; // @[TCU.scala 142:16]
  assign acc_io_input_bits_21 = router_io_acc_input_bits_21; // @[TCU.scala 142:16]
  assign acc_io_input_bits_22 = router_io_acc_input_bits_22; // @[TCU.scala 142:16]
  assign acc_io_input_bits_23 = router_io_acc_input_bits_23; // @[TCU.scala 142:16]
  assign acc_io_input_bits_24 = router_io_acc_input_bits_24; // @[TCU.scala 142:16]
  assign acc_io_input_bits_25 = router_io_acc_input_bits_25; // @[TCU.scala 142:16]
  assign acc_io_input_bits_26 = router_io_acc_input_bits_26; // @[TCU.scala 142:16]
  assign acc_io_input_bits_27 = router_io_acc_input_bits_27; // @[TCU.scala 142:16]
  assign acc_io_input_bits_28 = router_io_acc_input_bits_28; // @[TCU.scala 142:16]
  assign acc_io_input_bits_29 = router_io_acc_input_bits_29; // @[TCU.scala 142:16]
  assign acc_io_input_bits_30 = router_io_acc_input_bits_30; // @[TCU.scala 142:16]
  assign acc_io_input_bits_31 = router_io_acc_input_bits_31; // @[TCU.scala 142:16]
  assign acc_io_output_ready = router_io_acc_output_ready; // @[TCU.scala 143:24]
  assign acc_io_control_valid = acc_io_control_q_io_deq_valid; // @[TCU.scala 110:18]
  assign acc_io_control_bits_instruction_op = acc_io_control_q_io_deq_bits_instruction_op; // @[TCU.scala 110:18]
  assign acc_io_control_bits_instruction_sourceLeft = acc_io_control_q_io_deq_bits_instruction_sourceLeft; // @[TCU.scala 110:18]
  assign acc_io_control_bits_instruction_sourceRight = acc_io_control_q_io_deq_bits_instruction_sourceRight; // @[TCU.scala 110:18]
  assign acc_io_control_bits_instruction_dest = acc_io_control_q_io_deq_bits_instruction_dest; // @[TCU.scala 110:18]
  assign acc_io_control_bits_readAddress = acc_io_control_q_io_deq_bits_readAddress; // @[TCU.scala 110:18]
  assign acc_io_control_bits_writeAddress = acc_io_control_q_io_deq_bits_writeAddress; // @[TCU.scala 110:18]
  assign acc_io_control_bits_accumulate = acc_io_control_q_io_deq_bits_accumulate; // @[TCU.scala 110:18]
  assign acc_io_control_bits_write = acc_io_control_q_io_deq_bits_write; // @[TCU.scala 110:18]
  assign acc_io_control_bits_read = acc_io_control_q_io_deq_bits_read; // @[TCU.scala 110:18]
  assign acc_io_tracepoint = decoder_io_tracepoint; // @[TCU.scala 111:21]
  assign acc_io_programCounter = decoder_io_programCounter; // @[TCU.scala 112:25]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_portA_control_valid = decoder_io_memPortA_valid; // @[TCU.scala 124:17]
  assign mem_io_portA_control_bits_write = decoder_io_memPortA_bits_write; // @[TCU.scala 124:17]
  assign mem_io_portA_control_bits_address = decoder_io_memPortA_bits_address; // @[TCU.scala 124:17]
  assign mem_io_portA_input_valid = router_io_mem_input_valid; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_0 = router_io_mem_input_bits_0; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_1 = router_io_mem_input_bits_1; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_2 = router_io_mem_input_bits_2; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_3 = router_io_mem_input_bits_3; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_4 = router_io_mem_input_bits_4; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_5 = router_io_mem_input_bits_5; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_6 = router_io_mem_input_bits_6; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_7 = router_io_mem_input_bits_7; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_8 = router_io_mem_input_bits_8; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_9 = router_io_mem_input_bits_9; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_10 = router_io_mem_input_bits_10; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_11 = router_io_mem_input_bits_11; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_12 = router_io_mem_input_bits_12; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_13 = router_io_mem_input_bits_13; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_14 = router_io_mem_input_bits_14; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_15 = router_io_mem_input_bits_15; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_16 = router_io_mem_input_bits_16; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_17 = router_io_mem_input_bits_17; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_18 = router_io_mem_input_bits_18; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_19 = router_io_mem_input_bits_19; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_20 = router_io_mem_input_bits_20; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_21 = router_io_mem_input_bits_21; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_22 = router_io_mem_input_bits_22; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_23 = router_io_mem_input_bits_23; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_24 = router_io_mem_input_bits_24; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_25 = router_io_mem_input_bits_25; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_26 = router_io_mem_input_bits_26; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_27 = router_io_mem_input_bits_27; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_28 = router_io_mem_input_bits_28; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_29 = router_io_mem_input_bits_29; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_30 = router_io_mem_input_bits_30; // @[TCU.scala 136:15]
  assign mem_io_portA_input_bits_31 = router_io_mem_input_bits_31; // @[TCU.scala 136:15]
  assign mem_io_portA_output_ready = router_io_mem_output_ready; // @[TCU.scala 135:24]
  assign mem_io_portB_control_valid = decoder_io_memPortB_valid; // @[TCU.scala 148:17]
  assign mem_io_portB_control_bits_write = decoder_io_memPortB_bits_write; // @[TCU.scala 148:17]
  assign mem_io_portB_control_bits_address = decoder_io_memPortB_bits_address; // @[TCU.scala 148:17]
  assign mem_io_portB_input_valid = hostRouter_io_mem_input_valid; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_0 = hostRouter_io_mem_input_bits_0; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_1 = hostRouter_io_mem_input_bits_1; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_2 = hostRouter_io_mem_input_bits_2; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_3 = hostRouter_io_mem_input_bits_3; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_4 = hostRouter_io_mem_input_bits_4; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_5 = hostRouter_io_mem_input_bits_5; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_6 = hostRouter_io_mem_input_bits_6; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_7 = hostRouter_io_mem_input_bits_7; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_8 = hostRouter_io_mem_input_bits_8; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_9 = hostRouter_io_mem_input_bits_9; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_10 = hostRouter_io_mem_input_bits_10; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_11 = hostRouter_io_mem_input_bits_11; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_12 = hostRouter_io_mem_input_bits_12; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_13 = hostRouter_io_mem_input_bits_13; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_14 = hostRouter_io_mem_input_bits_14; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_15 = hostRouter_io_mem_input_bits_15; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_16 = hostRouter_io_mem_input_bits_16; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_17 = hostRouter_io_mem_input_bits_17; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_18 = hostRouter_io_mem_input_bits_18; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_19 = hostRouter_io_mem_input_bits_19; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_20 = hostRouter_io_mem_input_bits_20; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_21 = hostRouter_io_mem_input_bits_21; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_22 = hostRouter_io_mem_input_bits_22; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_23 = hostRouter_io_mem_input_bits_23; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_24 = hostRouter_io_mem_input_bits_24; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_25 = hostRouter_io_mem_input_bits_25; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_26 = hostRouter_io_mem_input_bits_26; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_27 = hostRouter_io_mem_input_bits_27; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_28 = hostRouter_io_mem_input_bits_28; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_29 = hostRouter_io_mem_input_bits_29; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_30 = hostRouter_io_mem_input_bits_30; // @[TCU.scala 149:15]
  assign mem_io_portB_input_bits_31 = hostRouter_io_mem_input_bits_31; // @[TCU.scala 149:15]
  assign mem_io_portB_output_ready = hostRouter_io_mem_output_ready; // @[TCU.scala 150:28]
  assign mem_io_tracepoint = decoder_io_tracepoint; // @[TCU.scala 122:21]
  assign mem_io_programCounter = decoder_io_programCounter; // @[TCU.scala 123:25]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_control_valid = decoder_io_dataflow_valid; // @[TCU.scala 133:21]
  assign router_io_control_bits_kind = decoder_io_dataflow_bits_kind; // @[TCU.scala 133:21]
  assign router_io_control_bits_size = decoder_io_dataflow_bits_size; // @[TCU.scala 133:21]
  assign router_io_mem_output_valid = mem_io_portA_output_valid; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_0 = mem_io_portA_output_bits_0; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_1 = mem_io_portA_output_bits_1; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_2 = mem_io_portA_output_bits_2; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_3 = mem_io_portA_output_bits_3; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_4 = mem_io_portA_output_bits_4; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_5 = mem_io_portA_output_bits_5; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_6 = mem_io_portA_output_bits_6; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_7 = mem_io_portA_output_bits_7; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_8 = mem_io_portA_output_bits_8; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_9 = mem_io_portA_output_bits_9; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_10 = mem_io_portA_output_bits_10; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_11 = mem_io_portA_output_bits_11; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_12 = mem_io_portA_output_bits_12; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_13 = mem_io_portA_output_bits_13; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_14 = mem_io_portA_output_bits_14; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_15 = mem_io_portA_output_bits_15; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_16 = mem_io_portA_output_bits_16; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_17 = mem_io_portA_output_bits_17; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_18 = mem_io_portA_output_bits_18; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_19 = mem_io_portA_output_bits_19; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_20 = mem_io_portA_output_bits_20; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_21 = mem_io_portA_output_bits_21; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_22 = mem_io_portA_output_bits_22; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_23 = mem_io_portA_output_bits_23; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_24 = mem_io_portA_output_bits_24; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_25 = mem_io_portA_output_bits_25; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_26 = mem_io_portA_output_bits_26; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_27 = mem_io_portA_output_bits_27; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_28 = mem_io_portA_output_bits_28; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_29 = mem_io_portA_output_bits_29; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_30 = mem_io_portA_output_bits_30; // @[TCU.scala 135:24]
  assign router_io_mem_output_bits_31 = mem_io_portA_output_bits_31; // @[TCU.scala 135:24]
  assign router_io_mem_input_ready = mem_io_portA_input_ready; // @[TCU.scala 136:15]
  assign router_io_array_input_ready = array_io_input_ready; // @[TCU.scala 138:18]
  assign router_io_array_output_valid = array_io_output_valid; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_0 = array_io_output_bits_0; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_1 = array_io_output_bits_1; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_2 = array_io_output_bits_2; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_3 = array_io_output_bits_3; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_4 = array_io_output_bits_4; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_5 = array_io_output_bits_5; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_6 = array_io_output_bits_6; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_7 = array_io_output_bits_7; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_8 = array_io_output_bits_8; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_9 = array_io_output_bits_9; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_10 = array_io_output_bits_10; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_11 = array_io_output_bits_11; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_12 = array_io_output_bits_12; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_13 = array_io_output_bits_13; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_14 = array_io_output_bits_14; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_15 = array_io_output_bits_15; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_16 = array_io_output_bits_16; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_17 = array_io_output_bits_17; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_18 = array_io_output_bits_18; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_19 = array_io_output_bits_19; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_20 = array_io_output_bits_20; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_21 = array_io_output_bits_21; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_22 = array_io_output_bits_22; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_23 = array_io_output_bits_23; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_24 = array_io_output_bits_24; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_25 = array_io_output_bits_25; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_26 = array_io_output_bits_26; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_27 = array_io_output_bits_27; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_28 = array_io_output_bits_28; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_29 = array_io_output_bits_29; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_30 = array_io_output_bits_30; // @[TCU.scala 139:26]
  assign router_io_array_output_bits_31 = array_io_output_bits_31; // @[TCU.scala 139:26]
  assign router_io_array_weightInput_ready = array_io_weight_ready; // @[TCU.scala 140:19]
  assign router_io_acc_output_valid = acc_io_output_valid; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_0 = acc_io_output_bits_0; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_1 = acc_io_output_bits_1; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_2 = acc_io_output_bits_2; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_3 = acc_io_output_bits_3; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_4 = acc_io_output_bits_4; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_5 = acc_io_output_bits_5; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_6 = acc_io_output_bits_6; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_7 = acc_io_output_bits_7; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_8 = acc_io_output_bits_8; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_9 = acc_io_output_bits_9; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_10 = acc_io_output_bits_10; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_11 = acc_io_output_bits_11; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_12 = acc_io_output_bits_12; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_13 = acc_io_output_bits_13; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_14 = acc_io_output_bits_14; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_15 = acc_io_output_bits_15; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_16 = acc_io_output_bits_16; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_17 = acc_io_output_bits_17; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_18 = acc_io_output_bits_18; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_19 = acc_io_output_bits_19; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_20 = acc_io_output_bits_20; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_21 = acc_io_output_bits_21; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_22 = acc_io_output_bits_22; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_23 = acc_io_output_bits_23; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_24 = acc_io_output_bits_24; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_25 = acc_io_output_bits_25; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_26 = acc_io_output_bits_26; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_27 = acc_io_output_bits_27; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_28 = acc_io_output_bits_28; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_29 = acc_io_output_bits_29; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_30 = acc_io_output_bits_30; // @[TCU.scala 143:24]
  assign router_io_acc_output_bits_31 = acc_io_output_bits_31; // @[TCU.scala 143:24]
  assign router_io_acc_input_ready = acc_io_input_ready; // @[TCU.scala 142:16]
  assign router_io_timeout = decoder_io_timeout; // @[TCU.scala 129:21]
  assign router_io_tracepoint = decoder_io_tracepoint; // @[TCU.scala 130:24]
  assign router_io_programCounter = decoder_io_programCounter; // @[TCU.scala 131:28]
  assign hostRouter_io_control_valid = decoder_io_hostDataflow_valid; // @[TCU.scala 146:25]
  assign hostRouter_io_control_bits_kind = decoder_io_hostDataflow_bits_kind; // @[TCU.scala 146:25]
  assign hostRouter_io_dram0_dataIn_valid = io_dram0_dataIn_valid; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_0 = io_dram0_dataIn_bits_0; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_1 = io_dram0_dataIn_bits_1; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_2 = io_dram0_dataIn_bits_2; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_3 = io_dram0_dataIn_bits_3; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_4 = io_dram0_dataIn_bits_4; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_5 = io_dram0_dataIn_bits_5; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_6 = io_dram0_dataIn_bits_6; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_7 = io_dram0_dataIn_bits_7; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_8 = io_dram0_dataIn_bits_8; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_9 = io_dram0_dataIn_bits_9; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_10 = io_dram0_dataIn_bits_10; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_11 = io_dram0_dataIn_bits_11; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_12 = io_dram0_dataIn_bits_12; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_13 = io_dram0_dataIn_bits_13; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_14 = io_dram0_dataIn_bits_14; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_15 = io_dram0_dataIn_bits_15; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_16 = io_dram0_dataIn_bits_16; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_17 = io_dram0_dataIn_bits_17; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_18 = io_dram0_dataIn_bits_18; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_19 = io_dram0_dataIn_bits_19; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_20 = io_dram0_dataIn_bits_20; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_21 = io_dram0_dataIn_bits_21; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_22 = io_dram0_dataIn_bits_22; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_23 = io_dram0_dataIn_bits_23; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_24 = io_dram0_dataIn_bits_24; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_25 = io_dram0_dataIn_bits_25; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_26 = io_dram0_dataIn_bits_26; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_27 = io_dram0_dataIn_bits_27; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_28 = io_dram0_dataIn_bits_28; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_29 = io_dram0_dataIn_bits_29; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_30 = io_dram0_dataIn_bits_30; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataIn_bits_31 = io_dram0_dataIn_bits_31; // @[TCU.scala 155:30]
  assign hostRouter_io_dram0_dataOut_ready = io_dram0_dataOut_ready; // @[TCU.scala 156:20]
  assign hostRouter_io_dram1_dataIn_valid = io_dram1_dataIn_valid; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_0 = io_dram1_dataIn_bits_0; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_1 = io_dram1_dataIn_bits_1; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_2 = io_dram1_dataIn_bits_2; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_3 = io_dram1_dataIn_bits_3; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_4 = io_dram1_dataIn_bits_4; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_5 = io_dram1_dataIn_bits_5; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_6 = io_dram1_dataIn_bits_6; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_7 = io_dram1_dataIn_bits_7; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_8 = io_dram1_dataIn_bits_8; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_9 = io_dram1_dataIn_bits_9; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_10 = io_dram1_dataIn_bits_10; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_11 = io_dram1_dataIn_bits_11; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_12 = io_dram1_dataIn_bits_12; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_13 = io_dram1_dataIn_bits_13; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_14 = io_dram1_dataIn_bits_14; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_15 = io_dram1_dataIn_bits_15; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_16 = io_dram1_dataIn_bits_16; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_17 = io_dram1_dataIn_bits_17; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_18 = io_dram1_dataIn_bits_18; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_19 = io_dram1_dataIn_bits_19; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_20 = io_dram1_dataIn_bits_20; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_21 = io_dram1_dataIn_bits_21; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_22 = io_dram1_dataIn_bits_22; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_23 = io_dram1_dataIn_bits_23; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_24 = io_dram1_dataIn_bits_24; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_25 = io_dram1_dataIn_bits_25; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_26 = io_dram1_dataIn_bits_26; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_27 = io_dram1_dataIn_bits_27; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_28 = io_dram1_dataIn_bits_28; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_29 = io_dram1_dataIn_bits_29; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_30 = io_dram1_dataIn_bits_30; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataIn_bits_31 = io_dram1_dataIn_bits_31; // @[TCU.scala 158:30]
  assign hostRouter_io_dram1_dataOut_ready = io_dram1_dataOut_ready; // @[TCU.scala 159:20]
  assign hostRouter_io_mem_output_valid = mem_io_portB_output_valid; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_0 = mem_io_portB_output_bits_0; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_1 = mem_io_portB_output_bits_1; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_2 = mem_io_portB_output_bits_2; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_3 = mem_io_portB_output_bits_3; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_4 = mem_io_portB_output_bits_4; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_5 = mem_io_portB_output_bits_5; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_6 = mem_io_portB_output_bits_6; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_7 = mem_io_portB_output_bits_7; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_8 = mem_io_portB_output_bits_8; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_9 = mem_io_portB_output_bits_9; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_10 = mem_io_portB_output_bits_10; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_11 = mem_io_portB_output_bits_11; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_12 = mem_io_portB_output_bits_12; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_13 = mem_io_portB_output_bits_13; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_14 = mem_io_portB_output_bits_14; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_15 = mem_io_portB_output_bits_15; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_16 = mem_io_portB_output_bits_16; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_17 = mem_io_portB_output_bits_17; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_18 = mem_io_portB_output_bits_18; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_19 = mem_io_portB_output_bits_19; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_20 = mem_io_portB_output_bits_20; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_21 = mem_io_portB_output_bits_21; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_22 = mem_io_portB_output_bits_22; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_23 = mem_io_portB_output_bits_23; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_24 = mem_io_portB_output_bits_24; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_25 = mem_io_portB_output_bits_25; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_26 = mem_io_portB_output_bits_26; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_27 = mem_io_portB_output_bits_27; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_28 = mem_io_portB_output_bits_28; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_29 = mem_io_portB_output_bits_29; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_30 = mem_io_portB_output_bits_30; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_output_bits_31 = mem_io_portB_output_bits_31; // @[TCU.scala 150:28]
  assign hostRouter_io_mem_input_ready = mem_io_portB_input_ready; // @[TCU.scala 149:15]
  assign acc_io_control_q_clock = clock;
  assign acc_io_control_q_reset = reset;
  assign acc_io_control_q_io_enq_valid = decoder_io_acc_valid; // @[TCU.scala 110:39]
  assign acc_io_control_q_io_enq_bits_instruction_op = decoder_io_acc_bits_instruction_op; // @[TCU.scala 110:39]
  assign acc_io_control_q_io_enq_bits_instruction_sourceLeft = decoder_io_acc_bits_instruction_sourceLeft; // @[TCU.scala 110:39]
  assign acc_io_control_q_io_enq_bits_instruction_sourceRight = decoder_io_acc_bits_instruction_sourceRight; // @[TCU.scala 110:39]
  assign acc_io_control_q_io_enq_bits_instruction_dest = decoder_io_acc_bits_instruction_dest; // @[TCU.scala 110:39]
  assign acc_io_control_q_io_enq_bits_readAddress = decoder_io_acc_bits_readAddress; // @[TCU.scala 110:39]
  assign acc_io_control_q_io_enq_bits_writeAddress = decoder_io_acc_bits_writeAddress; // @[TCU.scala 110:39]
  assign acc_io_control_q_io_enq_bits_accumulate = decoder_io_acc_bits_accumulate; // @[TCU.scala 110:39]
  assign acc_io_control_q_io_enq_bits_write = decoder_io_acc_bits_write; // @[TCU.scala 110:39]
  assign acc_io_control_q_io_enq_bits_read = decoder_io_acc_bits_read; // @[TCU.scala 110:39]
  assign acc_io_control_q_io_deq_ready = acc_io_control_ready; // @[TCU.scala 110:18]
  assign array_io_control_q_clock = clock;
  assign array_io_control_q_reset = reset;
  assign array_io_control_q_io_enq_valid = decoder_io_array_valid; // @[TCU.scala 117:41]
  assign array_io_control_q_io_enq_bits_load = decoder_io_array_bits_load; // @[TCU.scala 117:41]
  assign array_io_control_q_io_enq_bits_zeroes = decoder_io_array_bits_zeroes; // @[TCU.scala 117:41]
  assign array_io_control_q_io_deq_ready = array_io_control_ready; // @[TCU.scala 117:20]
endmodule
module Queue_30(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | ~full; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits = empty ? io_enq_bits : ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_32(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  ram [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | ~full; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits = empty ? io_enq_bits : ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram[initvar] = _RAND_0[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Counter_10(
  input        clock,
  input        reset,
  input        io_value_ready,
  output [7:0] io_value_bits,
  input        io_resetValue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] value; // @[Counter.scala 16:22]
  wire [7:0] _value_T_1 = value + 8'h1; // @[Counter.scala 24:22]
  assign io_value_bits = value; // @[Counter.scala 18:17]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 16:22]
      value <= 8'h0; // @[Counter.scala 16:22]
    end else if (io_resetValue) begin // @[Counter.scala 27:23]
      value <= 8'h0; // @[Counter.scala 28:11]
    end else if (io_value_ready) begin // @[Counter.scala 20:24]
      if (value == 8'hff) begin // @[Counter.scala 21:31]
        value <= 8'h0; // @[Counter.scala 22:13]
      end else begin
        value <= _value_T_1; // @[Counter.scala 24:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BurstSplitter(
  input          clock,
  input          reset,
  output         io_control_ready,
  input          io_control_valid,
  input  [7:0]   io_control_bits,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits_data,
  input          io_out_ready,
  output         io_out_valid,
  output [127:0] io_out_bits_data,
  output         io_out_bits_last
);
  wire  counter_clock; // @[Counter.scala 34:19]
  wire  counter_reset; // @[Counter.scala 34:19]
  wire  counter_io_value_ready; // @[Counter.scala 34:19]
  wire [7:0] counter_io_value_bits; // @[Counter.scala 34:19]
  wire  counter_io_resetValue; // @[Counter.scala 34:19]
  wire  _counter_io_resetValue_T = io_out_ready & io_out_valid; // @[Decoupled.scala 50:35]
  Counter_10 counter ( // @[Counter.scala 34:19]
    .clock(counter_clock),
    .reset(counter_reset),
    .io_value_ready(counter_io_value_ready),
    .io_value_bits(counter_io_value_bits),
    .io_resetValue(counter_io_resetValue)
  );
  assign io_control_ready = counter_io_value_bits == io_control_bits & _counter_io_resetValue_T; // @[MemBoundarySplitter.scala 45:51 48:22 52:22]
  assign io_in_ready = io_control_valid & io_out_ready; // @[MemBoundarySplitter.scala 41:35]
  assign io_out_valid = io_control_valid & io_in_valid; // @[MemBoundarySplitter.scala 40:36]
  assign io_out_bits_data = io_in_bits_data; // @[MemBoundarySplitter.scala 34:34]
  assign io_out_bits_last = counter_io_value_bits == io_control_bits; // @[MemBoundarySplitter.scala 45:30]
  assign counter_clock = clock;
  assign counter_reset = reset;
  assign counter_io_value_ready = counter_io_value_bits == io_control_bits ? 1'h0 : _counter_io_resetValue_T; // @[Counter.scala 36:22 MemBoundarySplitter.scala 45:51 51:28]
  assign counter_io_resetValue = counter_io_value_bits == io_control_bits & _counter_io_resetValue_T; // @[Counter.scala 35:21 MemBoundarySplitter.scala 45:51 47:27]
endmodule
module BurstSplitter_1(
  input          clock,
  input          reset,
  output         io_control_ready,
  input          io_control_valid,
  input  [7:0]   io_control_bits,
  output         io_in_ready,
  input          io_in_valid,
  input  [5:0]   io_in_bits_id,
  input  [127:0] io_in_bits_data,
  input  [15:0]  io_in_bits_strb,
  input          io_out_ready,
  output         io_out_valid,
  output [5:0]   io_out_bits_id,
  output [127:0] io_out_bits_data,
  output [15:0]  io_out_bits_strb,
  output         io_out_bits_last
);
  wire  counter_clock; // @[Counter.scala 34:19]
  wire  counter_reset; // @[Counter.scala 34:19]
  wire  counter_io_value_ready; // @[Counter.scala 34:19]
  wire [7:0] counter_io_value_bits; // @[Counter.scala 34:19]
  wire  counter_io_resetValue; // @[Counter.scala 34:19]
  wire  _counter_io_resetValue_T = io_out_ready & io_out_valid; // @[Decoupled.scala 50:35]
  Counter_10 counter ( // @[Counter.scala 34:19]
    .clock(counter_clock),
    .reset(counter_reset),
    .io_value_ready(counter_io_value_ready),
    .io_value_bits(counter_io_value_bits),
    .io_resetValue(counter_io_resetValue)
  );
  assign io_control_ready = counter_io_value_bits == io_control_bits & _counter_io_resetValue_T; // @[MemBoundarySplitter.scala 45:51 48:22 52:22]
  assign io_in_ready = io_control_valid & io_out_ready; // @[MemBoundarySplitter.scala 41:35]
  assign io_out_valid = io_control_valid & io_in_valid; // @[MemBoundarySplitter.scala 40:36]
  assign io_out_bits_id = io_in_bits_id; // @[MemBoundarySplitter.scala 34:34]
  assign io_out_bits_data = io_in_bits_data; // @[MemBoundarySplitter.scala 34:34]
  assign io_out_bits_strb = io_in_bits_strb; // @[MemBoundarySplitter.scala 34:34]
  assign io_out_bits_last = counter_io_value_bits == io_control_bits; // @[MemBoundarySplitter.scala 45:30]
  assign counter_clock = clock;
  assign counter_reset = reset;
  assign counter_io_value_ready = counter_io_value_bits == io_control_bits ? 1'h0 : _counter_io_resetValue_T; // @[Counter.scala 36:22 MemBoundarySplitter.scala 45:51 51:28]
  assign counter_io_resetValue = counter_io_value_bits == io_control_bits & _counter_io_resetValue_T; // @[Counter.scala 35:21 MemBoundarySplitter.scala 45:51 47:27]
endmodule
module Filter(
  output  io_control_ready,
  input   io_control_valid,
  input   io_control_bits,
  output  io_in_ready,
  input   io_in_valid,
  input   io_out_ready,
  output  io_out_valid
);
  assign io_control_ready = io_control_bits ? io_in_valid & io_out_ready : io_in_valid; // @[MemBoundarySplitter.scala 71:25 74:22 78:22]
  assign io_in_ready = io_control_bits ? io_control_valid & io_out_ready : io_control_valid; // @[MemBoundarySplitter.scala 71:25 73:17 77:17]
  assign io_out_valid = io_control_bits & (io_control_valid & io_in_valid); // @[MemBoundarySplitter.scala 71:25 72:18 76:18]
endmodule
module MemBoundarySplitter(
  input          clock,
  input          reset,
  output         io_in_writeAddress_ready,
  input          io_in_writeAddress_valid,
  input  [5:0]   io_in_writeAddress_bits_id,
  input  [31:0]  io_in_writeAddress_bits_addr,
  input  [7:0]   io_in_writeAddress_bits_len,
  input  [2:0]   io_in_writeAddress_bits_size,
  input  [1:0]   io_in_writeAddress_bits_burst,
  input  [1:0]   io_in_writeAddress_bits_lock,
  input  [3:0]   io_in_writeAddress_bits_cache,
  input  [2:0]   io_in_writeAddress_bits_prot,
  input  [3:0]   io_in_writeAddress_bits_qos,
  output         io_in_writeData_ready,
  input          io_in_writeData_valid,
  input  [5:0]   io_in_writeData_bits_id,
  input  [127:0] io_in_writeData_bits_data,
  input  [15:0]  io_in_writeData_bits_strb,
  input          io_in_writeResponse_ready,
  output         io_in_writeResponse_valid,
  output         io_in_readAddress_ready,
  input          io_in_readAddress_valid,
  input  [5:0]   io_in_readAddress_bits_id,
  input  [31:0]  io_in_readAddress_bits_addr,
  input  [7:0]   io_in_readAddress_bits_len,
  input  [2:0]   io_in_readAddress_bits_size,
  input  [1:0]   io_in_readAddress_bits_burst,
  input  [1:0]   io_in_readAddress_bits_lock,
  input  [3:0]   io_in_readAddress_bits_cache,
  input  [2:0]   io_in_readAddress_bits_prot,
  input  [3:0]   io_in_readAddress_bits_qos,
  input          io_in_readData_ready,
  output         io_in_readData_valid,
  output [127:0] io_in_readData_bits_data,
  output         io_in_readData_bits_last,
  input          io_out_writeAddress_ready,
  output         io_out_writeAddress_valid,
  output [5:0]   io_out_writeAddress_bits_id,
  output [31:0]  io_out_writeAddress_bits_addr,
  output [7:0]   io_out_writeAddress_bits_len,
  output [2:0]   io_out_writeAddress_bits_size,
  output [1:0]   io_out_writeAddress_bits_burst,
  output [1:0]   io_out_writeAddress_bits_lock,
  output [3:0]   io_out_writeAddress_bits_cache,
  output [2:0]   io_out_writeAddress_bits_prot,
  output [3:0]   io_out_writeAddress_bits_qos,
  input          io_out_writeData_ready,
  output         io_out_writeData_valid,
  output [5:0]   io_out_writeData_bits_id,
  output [127:0] io_out_writeData_bits_data,
  output [15:0]  io_out_writeData_bits_strb,
  output         io_out_writeData_bits_last,
  output         io_out_writeResponse_ready,
  input          io_out_writeResponse_valid,
  input          io_out_readAddress_ready,
  output         io_out_readAddress_valid,
  output [5:0]   io_out_readAddress_bits_id,
  output [31:0]  io_out_readAddress_bits_addr,
  output [7:0]   io_out_readAddress_bits_len,
  output [2:0]   io_out_readAddress_bits_size,
  output [1:0]   io_out_readAddress_bits_burst,
  output [1:0]   io_out_readAddress_bits_lock,
  output [3:0]   io_out_readAddress_bits_cache,
  output [2:0]   io_out_readAddress_bits_prot,
  output [3:0]   io_out_readAddress_bits_qos,
  output         io_out_readData_ready,
  input          io_out_readData_valid,
  input  [127:0] io_out_readData_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  readDataQueue_clock; // @[MemBoundarySplitter.scala 111:29]
  wire  readDataQueue_reset; // @[MemBoundarySplitter.scala 111:29]
  wire  readDataQueue_io_enq_ready; // @[MemBoundarySplitter.scala 111:29]
  wire  readDataQueue_io_enq_valid; // @[MemBoundarySplitter.scala 111:29]
  wire [7:0] readDataQueue_io_enq_bits; // @[MemBoundarySplitter.scala 111:29]
  wire  readDataQueue_io_deq_ready; // @[MemBoundarySplitter.scala 111:29]
  wire  readDataQueue_io_deq_valid; // @[MemBoundarySplitter.scala 111:29]
  wire [7:0] readDataQueue_io_deq_bits; // @[MemBoundarySplitter.scala 111:29]
  wire  writeDataQueue_clock; // @[MemBoundarySplitter.scala 114:30]
  wire  writeDataQueue_reset; // @[MemBoundarySplitter.scala 114:30]
  wire  writeDataQueue_io_enq_ready; // @[MemBoundarySplitter.scala 114:30]
  wire  writeDataQueue_io_enq_valid; // @[MemBoundarySplitter.scala 114:30]
  wire [7:0] writeDataQueue_io_enq_bits; // @[MemBoundarySplitter.scala 114:30]
  wire  writeDataQueue_io_deq_ready; // @[MemBoundarySplitter.scala 114:30]
  wire  writeDataQueue_io_deq_valid; // @[MemBoundarySplitter.scala 114:30]
  wire [7:0] writeDataQueue_io_deq_bits; // @[MemBoundarySplitter.scala 114:30]
  wire  writeResponseQueue_clock; // @[MemBoundarySplitter.scala 117:34]
  wire  writeResponseQueue_reset; // @[MemBoundarySplitter.scala 117:34]
  wire  writeResponseQueue_io_enq_ready; // @[MemBoundarySplitter.scala 117:34]
  wire  writeResponseQueue_io_enq_valid; // @[MemBoundarySplitter.scala 117:34]
  wire  writeResponseQueue_io_enq_bits; // @[MemBoundarySplitter.scala 117:34]
  wire  writeResponseQueue_io_deq_ready; // @[MemBoundarySplitter.scala 117:34]
  wire  writeResponseQueue_io_deq_valid; // @[MemBoundarySplitter.scala 117:34]
  wire  writeResponseQueue_io_deq_bits; // @[MemBoundarySplitter.scala 117:34]
  wire  readMerger_clock; // @[MemBoundarySplitter.scala 121:26]
  wire  readMerger_reset; // @[MemBoundarySplitter.scala 121:26]
  wire  readMerger_io_control_ready; // @[MemBoundarySplitter.scala 121:26]
  wire  readMerger_io_control_valid; // @[MemBoundarySplitter.scala 121:26]
  wire [7:0] readMerger_io_control_bits; // @[MemBoundarySplitter.scala 121:26]
  wire  readMerger_io_in_ready; // @[MemBoundarySplitter.scala 121:26]
  wire  readMerger_io_in_valid; // @[MemBoundarySplitter.scala 121:26]
  wire [127:0] readMerger_io_in_bits_data; // @[MemBoundarySplitter.scala 121:26]
  wire  readMerger_io_out_ready; // @[MemBoundarySplitter.scala 121:26]
  wire  readMerger_io_out_valid; // @[MemBoundarySplitter.scala 121:26]
  wire [127:0] readMerger_io_out_bits_data; // @[MemBoundarySplitter.scala 121:26]
  wire  readMerger_io_out_bits_last; // @[MemBoundarySplitter.scala 121:26]
  wire  writeSplitter_clock; // @[MemBoundarySplitter.scala 125:29]
  wire  writeSplitter_reset; // @[MemBoundarySplitter.scala 125:29]
  wire  writeSplitter_io_control_ready; // @[MemBoundarySplitter.scala 125:29]
  wire  writeSplitter_io_control_valid; // @[MemBoundarySplitter.scala 125:29]
  wire [7:0] writeSplitter_io_control_bits; // @[MemBoundarySplitter.scala 125:29]
  wire  writeSplitter_io_in_ready; // @[MemBoundarySplitter.scala 125:29]
  wire  writeSplitter_io_in_valid; // @[MemBoundarySplitter.scala 125:29]
  wire [5:0] writeSplitter_io_in_bits_id; // @[MemBoundarySplitter.scala 125:29]
  wire [127:0] writeSplitter_io_in_bits_data; // @[MemBoundarySplitter.scala 125:29]
  wire [15:0] writeSplitter_io_in_bits_strb; // @[MemBoundarySplitter.scala 125:29]
  wire  writeSplitter_io_out_ready; // @[MemBoundarySplitter.scala 125:29]
  wire  writeSplitter_io_out_valid; // @[MemBoundarySplitter.scala 125:29]
  wire [5:0] writeSplitter_io_out_bits_id; // @[MemBoundarySplitter.scala 125:29]
  wire [127:0] writeSplitter_io_out_bits_data; // @[MemBoundarySplitter.scala 125:29]
  wire [15:0] writeSplitter_io_out_bits_strb; // @[MemBoundarySplitter.scala 125:29]
  wire  writeSplitter_io_out_bits_last; // @[MemBoundarySplitter.scala 125:29]
  wire  writeResponseFilter_io_control_ready; // @[MemBoundarySplitter.scala 129:35]
  wire  writeResponseFilter_io_control_valid; // @[MemBoundarySplitter.scala 129:35]
  wire  writeResponseFilter_io_control_bits; // @[MemBoundarySplitter.scala 129:35]
  wire  writeResponseFilter_io_in_ready; // @[MemBoundarySplitter.scala 129:35]
  wire  writeResponseFilter_io_in_valid; // @[MemBoundarySplitter.scala 129:35]
  wire  writeResponseFilter_io_out_ready; // @[MemBoundarySplitter.scala 129:35]
  wire  writeResponseFilter_io_out_valid; // @[MemBoundarySplitter.scala 129:35]
  wire  readEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  readEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_clock; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_reset; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_2_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueuer_io_out_2_valid; // @[MultiEnqueue.scala 182:43]
  reg [11:0] readAddressCounter; // @[MemBoundarySplitter.scala 137:35]
  reg [7:0] readLenCounter; // @[MemBoundarySplitter.scala 140:31]
  reg [11:0] writeAddressCounter; // @[MemBoundarySplitter.scala 141:36]
  reg [7:0] writeLenCounter; // @[MemBoundarySplitter.scala 144:32]
  wire [12:0] lengthBytes = io_in_readAddress_bits_len * 5'h10; // @[MemBoundarySplitter.scala 105:30]
  wire [31:0] _GEN_141 = io_in_readAddress_bits_addr % 32'h1000; // @[MemBoundarySplitter.scala 106:45]
  wire [12:0] _T_3 = 13'h1001 - lengthBytes; // @[MemBoundarySplitter.scala 106:79]
  wire  _T_5 = lengthBytes > 13'h1000 | _GEN_141[12:0] > _T_3; // @[MemBoundarySplitter.scala 106:32]
  wire [31:0] _GEN_125 = {{20'd0}, readAddressCounter}; // @[MemBoundarySplitter.scala 151:44]
  wire [31:0] addr = io_in_readAddress_bits_addr + _GEN_125; // @[MemBoundarySplitter.scala 151:44]
  wire [31:0] _GEN_142 = addr % 32'h1000; // @[MemBoundarySplitter.scala 153:27]
  wire [12:0] availableAddresses = 13'h1000 - _GEN_142[12:0]; // @[MemBoundarySplitter.scala 153:19]
  wire [12:0] availableBeats = availableAddresses / 5'h10; // @[MemBoundarySplitter.scala 154:45]
  wire  _len_T = readLenCounter == 8'h0; // @[MemBoundarySplitter.scala 156:22]
  wire [12:0] _GEN_126 = {{5'd0}, readLenCounter}; // @[MemBoundarySplitter.scala 109:43]
  wire [12:0] _len_T_2 = availableBeats > _GEN_126 ? {{5'd0}, readLenCounter} : availableBeats; // @[MemBoundarySplitter.scala 109:40]
  wire [12:0] _len_T_3 = _len_T ? availableBeats : _len_T_2; // @[MemBoundarySplitter.scala 155:18]
  wire [12:0] len = _len_T_3 - 13'h1; // @[MemBoundarySplitter.scala 159:7]
  wire [12:0] _GEN_127 = {{5'd0}, io_in_readAddress_bits_len}; // @[MemBoundarySplitter.scala 182:54]
  wire [12:0] _readLenCounter_T_1 = _GEN_127 - len; // @[MemBoundarySplitter.scala 182:54]
  wire [12:0] _GEN_0 = io_in_readAddress_valid & readEnqueuer_io_in_ready ? availableAddresses : {{1'd0},
    readAddressCounter}; // @[MemBoundarySplitter.scala 180:46 181:28 137:35]
  wire [12:0] _GEN_1 = io_in_readAddress_valid & readEnqueuer_io_in_ready ? _readLenCounter_T_1 : {{5'd0},
    readLenCounter}; // @[MemBoundarySplitter.scala 180:46 182:24 140:31]
  wire  _T_9 = io_out_readAddress_ready & io_out_readAddress_valid; // @[Decoupled.scala 50:35]
  wire [11:0] _GEN_2 = _T_9 ? 12'h0 : readAddressCounter; // @[MemBoundarySplitter.scala 193:37 194:28 137:35]
  wire [7:0] _GEN_3 = _T_9 ? 8'h0 : readLenCounter; // @[MemBoundarySplitter.scala 193:37 195:24 140:31]
  wire [12:0] _GEN_129 = {{1'd0}, readAddressCounter}; // @[MemBoundarySplitter.scala 208:50]
  wire [12:0] _readAddressCounter_T_1 = _GEN_129 + availableAddresses; // @[MemBoundarySplitter.scala 208:50]
  wire [12:0] _readLenCounter_T_3 = len + 13'h1; // @[MemBoundarySplitter.scala 210:49]
  wire [12:0] _readLenCounter_T_5 = _GEN_126 - _readLenCounter_T_3; // @[MemBoundarySplitter.scala 210:42]
  wire [12:0] _GEN_4 = _T_9 ? _readAddressCounter_T_1 : {{1'd0}, readAddressCounter}; // @[MemBoundarySplitter.scala 206:37 208:28 137:35]
  wire [12:0] _GEN_5 = _T_9 ? _readLenCounter_T_5 : {{5'd0}, readLenCounter}; // @[MemBoundarySplitter.scala 206:37 210:24 140:31]
  wire  _GEN_7 = _GEN_126 <= availableBeats & io_out_readAddress_ready; // @[MemBoundarySplitter.scala 184:50 187:31 Decoupled.scala 88:20]
  wire [7:0] address_len = len[7:0]; // @[MemBoundarySplitter.scala 161:23 168:17]
  wire [12:0] _GEN_18 = _GEN_126 <= availableBeats ? {{1'd0}, _GEN_2} : _GEN_4; // @[MemBoundarySplitter.scala 184:50]
  wire [12:0] _GEN_19 = _GEN_126 <= availableBeats ? {{5'd0}, _GEN_3} : _GEN_5; // @[MemBoundarySplitter.scala 184:50]
  wire  _GEN_20 = _len_T & io_in_readAddress_valid; // @[MemBoundarySplitter.scala 170:34 MultiEnqueue.scala 84:17]
  wire  _GEN_21 = _len_T & io_out_readAddress_ready; // @[MemBoundarySplitter.scala 170:34 ReadyValid.scala 19:11]
  wire  ready_io_out_readAddress_w_valid = readEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_22 = _len_T ? ready_io_out_readAddress_w_valid : io_in_readAddress_valid; // @[MemBoundarySplitter.scala 170:34 MultiEnqueue.scala 85:10]
  wire  ready_readDataQueue_io_enq_w_ready = readDataQueue_io_enq_ready; // @[ReadyValid.scala 16:17 MultiEnqueue.scala 86:10]
  wire  _GEN_32 = _len_T & ready_readDataQueue_io_enq_w_ready; // @[MemBoundarySplitter.scala 170:34 ReadyValid.scala 19:11]
  wire  ready_readDataQueue_io_enq_w_valid = readEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_33 = _len_T & ready_readDataQueue_io_enq_w_valid; // @[MemBoundarySplitter.scala 170:34 MultiEnqueue.scala 86:10]
  wire  _GEN_35 = _len_T ? 1'h0 : _GEN_7; // @[MemBoundarySplitter.scala 170:34 Decoupled.scala 88:20]
  wire [12:0] _GEN_36 = _len_T ? _GEN_0 : _GEN_18; // @[MemBoundarySplitter.scala 170:34]
  wire [12:0] _GEN_37 = _len_T ? _GEN_1 : _GEN_19; // @[MemBoundarySplitter.scala 170:34]
  wire [12:0] _GEN_54 = _T_5 ? _GEN_36 : {{1'd0}, readAddressCounter}; // @[MemBoundarySplitter.scala 137:35 150:74]
  wire [12:0] _GEN_55 = _T_5 ? _GEN_37 : {{5'd0}, readLenCounter}; // @[MemBoundarySplitter.scala 140:31 150:74]
  wire [12:0] lengthBytes_1 = io_in_writeAddress_bits_len * 5'h10; // @[MemBoundarySplitter.scala 105:30]
  wire [31:0] _GEN_143 = io_in_writeAddress_bits_addr % 32'h1000; // @[MemBoundarySplitter.scala 106:45]
  wire [12:0] _T_14 = 13'h1001 - lengthBytes_1; // @[MemBoundarySplitter.scala 106:79]
  wire  _T_16 = lengthBytes_1 > 13'h1000 | _GEN_143[12:0] > _T_14; // @[MemBoundarySplitter.scala 106:32]
  wire [31:0] _GEN_131 = {{20'd0}, writeAddressCounter}; // @[MemBoundarySplitter.scala 225:45]
  wire [31:0] addr_1 = io_in_writeAddress_bits_addr + _GEN_131; // @[MemBoundarySplitter.scala 225:45]
  wire [31:0] _GEN_144 = addr_1 % 32'h1000; // @[MemBoundarySplitter.scala 227:27]
  wire [12:0] availableAddresses_1 = 13'h1000 - _GEN_144[12:0]; // @[MemBoundarySplitter.scala 227:19]
  wire [12:0] availableBeats_1 = availableAddresses_1 / 5'h10; // @[MemBoundarySplitter.scala 228:45]
  wire  _len_T_5 = writeLenCounter == 8'h0; // @[MemBoundarySplitter.scala 230:23]
  wire [12:0] _GEN_132 = {{5'd0}, writeLenCounter}; // @[MemBoundarySplitter.scala 109:43]
  wire [12:0] _len_T_7 = availableBeats_1 > _GEN_132 ? {{5'd0}, writeLenCounter} : availableBeats_1; // @[MemBoundarySplitter.scala 109:40]
  wire [12:0] _len_T_8 = _len_T_5 ? availableBeats_1 : _len_T_7; // @[MemBoundarySplitter.scala 229:18]
  wire [12:0] len_1 = _len_T_8 - 13'h1; // @[MemBoundarySplitter.scala 233:7]
  wire  _T_18 = io_in_writeAddress_valid & writeEnqueuer_io_in_ready; // @[MemBoundarySplitter.scala 256:37]
  wire [12:0] _GEN_133 = {{5'd0}, io_in_writeAddress_bits_len}; // @[MemBoundarySplitter.scala 258:56]
  wire [12:0] _writeLenCounter_T_1 = _GEN_133 - len_1; // @[MemBoundarySplitter.scala 258:56]
  wire [12:0] _GEN_56 = io_in_writeAddress_valid & writeEnqueuer_io_in_ready ? availableAddresses_1 : {{1'd0},
    writeAddressCounter}; // @[MemBoundarySplitter.scala 256:47 257:29 141:36]
  wire [12:0] _GEN_57 = io_in_writeAddress_valid & writeEnqueuer_io_in_ready ? _writeLenCounter_T_1 : {{5'd0},
    writeLenCounter}; // @[MemBoundarySplitter.scala 256:47 258:25 144:32]
  wire  _T_19 = _GEN_132 <= availableBeats_1; // @[MemBoundarySplitter.scala 260:32]
  wire [11:0] _GEN_58 = _T_18 ? 12'h0 : writeAddressCounter; // @[MemBoundarySplitter.scala 272:47 273:29 141:36]
  wire [7:0] _GEN_59 = _T_18 ? 8'h0 : writeLenCounter; // @[MemBoundarySplitter.scala 272:47 274:25 144:32]
  wire [12:0] _GEN_135 = {{1'd0}, writeAddressCounter}; // @[MemBoundarySplitter.scala 290:52]
  wire [12:0] _writeAddressCounter_T_1 = _GEN_135 + availableAddresses_1; // @[MemBoundarySplitter.scala 290:52]
  wire [12:0] _writeLenCounter_T_3 = len_1 + 13'h1; // @[MemBoundarySplitter.scala 292:51]
  wire [12:0] _writeLenCounter_T_5 = _GEN_132 - _writeLenCounter_T_3; // @[MemBoundarySplitter.scala 292:44]
  wire [12:0] _GEN_60 = _T_18 ? _writeAddressCounter_T_1 : {{1'd0}, writeAddressCounter}; // @[MemBoundarySplitter.scala 288:47 290:29 141:36]
  wire [12:0] _GEN_61 = _T_18 ? _writeLenCounter_T_5 : {{5'd0}, writeLenCounter}; // @[MemBoundarySplitter.scala 288:47 292:25 144:32]
  wire  ready_io_out_writeAddress_w_1_valid = writeEnqueuer_io_out_0_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_64 = _GEN_132 <= availableBeats_1 ? ready_io_out_writeAddress_w_1_valid :
    ready_io_out_writeAddress_w_1_valid; // @[MemBoundarySplitter.scala 260:51 MultiEnqueue.scala 115:{10,10}]
  wire [7:0] address_1_len = len_1[7:0]; // @[MemBoundarySplitter.scala 235:23 242:17]
  wire  ready_writeDataQueue_io_enq_w_1_ready = writeDataQueue_io_enq_ready; // @[MultiEnqueue.scala 116:10 ReadyValid.scala 16:17]
  wire  _GEN_74 = _GEN_132 <= availableBeats_1 ? ready_writeDataQueue_io_enq_w_1_ready :
    ready_writeDataQueue_io_enq_w_1_ready; // @[MemBoundarySplitter.scala 260:51 ReadyValid.scala 19:{11,11}]
  wire  ready_writeDataQueue_io_enq_w_1_valid = writeEnqueuer_io_out_1_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_75 = _GEN_132 <= availableBeats_1 ? ready_writeDataQueue_io_enq_w_1_valid :
    ready_writeDataQueue_io_enq_w_1_valid; // @[MemBoundarySplitter.scala 260:51 MultiEnqueue.scala 116:{10,10}]
  wire  ready_writeResponseQueue_io_enq_w_1_ready = writeResponseQueue_io_enq_ready; // @[MultiEnqueue.scala 117:10 ReadyValid.scala 16:17]
  wire  _GEN_77 = _GEN_132 <= availableBeats_1 ? ready_writeResponseQueue_io_enq_w_1_ready :
    ready_writeResponseQueue_io_enq_w_1_ready; // @[MemBoundarySplitter.scala 260:51 ReadyValid.scala 19:{11,11}]
  wire  ready_writeResponseQueue_io_enq_w_1_valid = writeEnqueuer_io_out_2_valid; // @[ReadyValid.scala 16:17 18:13]
  wire  _GEN_78 = _GEN_132 <= availableBeats_1 ? ready_writeResponseQueue_io_enq_w_1_valid :
    ready_writeResponseQueue_io_enq_w_1_valid; // @[MemBoundarySplitter.scala 260:51 MultiEnqueue.scala 117:{10,10}]
  wire  _GEN_80 = _GEN_132 <= availableBeats_1 & writeEnqueuer_io_in_ready; // @[MemBoundarySplitter.scala 260:51 271:32 Decoupled.scala 88:20]
  wire [12:0] _GEN_81 = _GEN_132 <= availableBeats_1 ? {{1'd0}, _GEN_58} : _GEN_60; // @[MemBoundarySplitter.scala 260:51]
  wire [12:0] _GEN_82 = _GEN_132 <= availableBeats_1 ? {{5'd0}, _GEN_59} : _GEN_61; // @[MemBoundarySplitter.scala 260:51]
  wire  _GEN_85 = _len_T_5 ? ready_io_out_writeAddress_w_1_valid : _GEN_64; // @[MemBoundarySplitter.scala 244:35 MultiEnqueue.scala 115:10]
  wire  _GEN_95 = _len_T_5 ? ready_writeDataQueue_io_enq_w_1_ready : _GEN_74; // @[MemBoundarySplitter.scala 244:35 ReadyValid.scala 19:11]
  wire  _GEN_96 = _len_T_5 ? ready_writeDataQueue_io_enq_w_1_valid : _GEN_75; // @[MemBoundarySplitter.scala 244:35 MultiEnqueue.scala 116:10]
  wire  _GEN_98 = _len_T_5 ? ready_writeResponseQueue_io_enq_w_1_ready : _GEN_77; // @[MemBoundarySplitter.scala 244:35 ReadyValid.scala 19:11]
  wire  _GEN_99 = _len_T_5 ? ready_writeResponseQueue_io_enq_w_1_valid : _GEN_78; // @[MemBoundarySplitter.scala 244:35 MultiEnqueue.scala 117:10]
  wire  _GEN_100 = _len_T_5 ? 1'h0 : _T_19; // @[MemBoundarySplitter.scala 244:35 MultiEnqueue.scala 117:10]
  wire  _GEN_101 = _len_T_5 ? 1'h0 : _GEN_80; // @[MemBoundarySplitter.scala 244:35 Decoupled.scala 88:20]
  wire [12:0] _GEN_102 = _len_T_5 ? _GEN_56 : _GEN_81; // @[MemBoundarySplitter.scala 244:35]
  wire [12:0] _GEN_103 = _len_T_5 ? _GEN_57 : _GEN_82; // @[MemBoundarySplitter.scala 244:35]
  wire [12:0] _GEN_123 = _T_16 ? _GEN_102 : {{1'd0}, writeAddressCounter}; // @[MemBoundarySplitter.scala 141:36 224:76]
  wire [12:0] _GEN_124 = _T_16 ? _GEN_103 : {{5'd0}, writeLenCounter}; // @[MemBoundarySplitter.scala 144:32 224:76]
  wire [12:0] _GEN_137 = reset ? 13'h0 : _GEN_54; // @[MemBoundarySplitter.scala 137:{35,35}]
  wire [12:0] _GEN_138 = reset ? 13'h0 : _GEN_55; // @[MemBoundarySplitter.scala 140:{31,31}]
  wire [12:0] _GEN_139 = reset ? 13'h0 : _GEN_123; // @[MemBoundarySplitter.scala 141:{36,36}]
  wire [12:0] _GEN_140 = reset ? 13'h0 : _GEN_124; // @[MemBoundarySplitter.scala 144:{32,32}]
  Queue_30 readDataQueue ( // @[MemBoundarySplitter.scala 111:29]
    .clock(readDataQueue_clock),
    .reset(readDataQueue_reset),
    .io_enq_ready(readDataQueue_io_enq_ready),
    .io_enq_valid(readDataQueue_io_enq_valid),
    .io_enq_bits(readDataQueue_io_enq_bits),
    .io_deq_ready(readDataQueue_io_deq_ready),
    .io_deq_valid(readDataQueue_io_deq_valid),
    .io_deq_bits(readDataQueue_io_deq_bits)
  );
  Queue_30 writeDataQueue ( // @[MemBoundarySplitter.scala 114:30]
    .clock(writeDataQueue_clock),
    .reset(writeDataQueue_reset),
    .io_enq_ready(writeDataQueue_io_enq_ready),
    .io_enq_valid(writeDataQueue_io_enq_valid),
    .io_enq_bits(writeDataQueue_io_enq_bits),
    .io_deq_ready(writeDataQueue_io_deq_ready),
    .io_deq_valid(writeDataQueue_io_deq_valid),
    .io_deq_bits(writeDataQueue_io_deq_bits)
  );
  Queue_32 writeResponseQueue ( // @[MemBoundarySplitter.scala 117:34]
    .clock(writeResponseQueue_clock),
    .reset(writeResponseQueue_reset),
    .io_enq_ready(writeResponseQueue_io_enq_ready),
    .io_enq_valid(writeResponseQueue_io_enq_valid),
    .io_enq_bits(writeResponseQueue_io_enq_bits),
    .io_deq_ready(writeResponseQueue_io_deq_ready),
    .io_deq_valid(writeResponseQueue_io_deq_valid),
    .io_deq_bits(writeResponseQueue_io_deq_bits)
  );
  BurstSplitter readMerger ( // @[MemBoundarySplitter.scala 121:26]
    .clock(readMerger_clock),
    .reset(readMerger_reset),
    .io_control_ready(readMerger_io_control_ready),
    .io_control_valid(readMerger_io_control_valid),
    .io_control_bits(readMerger_io_control_bits),
    .io_in_ready(readMerger_io_in_ready),
    .io_in_valid(readMerger_io_in_valid),
    .io_in_bits_data(readMerger_io_in_bits_data),
    .io_out_ready(readMerger_io_out_ready),
    .io_out_valid(readMerger_io_out_valid),
    .io_out_bits_data(readMerger_io_out_bits_data),
    .io_out_bits_last(readMerger_io_out_bits_last)
  );
  BurstSplitter_1 writeSplitter ( // @[MemBoundarySplitter.scala 125:29]
    .clock(writeSplitter_clock),
    .reset(writeSplitter_reset),
    .io_control_ready(writeSplitter_io_control_ready),
    .io_control_valid(writeSplitter_io_control_valid),
    .io_control_bits(writeSplitter_io_control_bits),
    .io_in_ready(writeSplitter_io_in_ready),
    .io_in_valid(writeSplitter_io_in_valid),
    .io_in_bits_id(writeSplitter_io_in_bits_id),
    .io_in_bits_data(writeSplitter_io_in_bits_data),
    .io_in_bits_strb(writeSplitter_io_in_bits_strb),
    .io_out_ready(writeSplitter_io_out_ready),
    .io_out_valid(writeSplitter_io_out_valid),
    .io_out_bits_id(writeSplitter_io_out_bits_id),
    .io_out_bits_data(writeSplitter_io_out_bits_data),
    .io_out_bits_strb(writeSplitter_io_out_bits_strb),
    .io_out_bits_last(writeSplitter_io_out_bits_last)
  );
  Filter writeResponseFilter ( // @[MemBoundarySplitter.scala 129:35]
    .io_control_ready(writeResponseFilter_io_control_ready),
    .io_control_valid(writeResponseFilter_io_control_valid),
    .io_control_bits(writeResponseFilter_io_control_bits),
    .io_in_ready(writeResponseFilter_io_in_ready),
    .io_in_valid(writeResponseFilter_io_in_valid),
    .io_out_ready(writeResponseFilter_io_out_ready),
    .io_out_valid(writeResponseFilter_io_out_valid)
  );
  MultiEnqueue_1 readEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(readEnqueuer_clock),
    .reset(readEnqueuer_reset),
    .io_in_ready(readEnqueuer_io_in_ready),
    .io_in_valid(readEnqueuer_io_in_valid),
    .io_out_0_ready(readEnqueuer_io_out_0_ready),
    .io_out_0_valid(readEnqueuer_io_out_0_valid),
    .io_out_1_ready(readEnqueuer_io_out_1_ready),
    .io_out_1_valid(readEnqueuer_io_out_1_valid)
  );
  MultiEnqueue_2 writeEnqueuer ( // @[MultiEnqueue.scala 182:43]
    .clock(writeEnqueuer_clock),
    .reset(writeEnqueuer_reset),
    .io_in_ready(writeEnqueuer_io_in_ready),
    .io_in_valid(writeEnqueuer_io_in_valid),
    .io_out_0_ready(writeEnqueuer_io_out_0_ready),
    .io_out_0_valid(writeEnqueuer_io_out_0_valid),
    .io_out_1_ready(writeEnqueuer_io_out_1_ready),
    .io_out_1_valid(writeEnqueuer_io_out_1_valid),
    .io_out_2_ready(writeEnqueuer_io_out_2_ready),
    .io_out_2_valid(writeEnqueuer_io_out_2_valid)
  );
  assign io_in_writeAddress_ready = _T_16 ? _GEN_101 : writeEnqueuer_io_in_ready; // @[MemBoundarySplitter.scala 224:76 296:30]
  assign io_in_writeData_ready = writeSplitter_io_in_ready; // @[MemBoundarySplitter.scala 127:23]
  assign io_in_writeResponse_valid = writeResponseFilter_io_out_valid; // @[MemBoundarySplitter.scala 132:23]
  assign io_in_readAddress_ready = _T_5 ? _GEN_35 : readEnqueuer_io_in_ready; // @[MemBoundarySplitter.scala 150:74 214:29]
  assign io_in_readData_valid = readMerger_io_out_valid; // @[MemBoundarySplitter.scala 124:18]
  assign io_in_readData_bits_data = readMerger_io_out_bits_data; // @[MemBoundarySplitter.scala 124:18]
  assign io_in_readData_bits_last = readMerger_io_out_bits_last; // @[MemBoundarySplitter.scala 124:18]
  assign io_out_writeAddress_valid = _T_16 ? _GEN_85 : ready_io_out_writeAddress_w_1_valid; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 115:10]
  assign io_out_writeAddress_bits_id = io_in_writeAddress_bits_id; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 115:10]
  assign io_out_writeAddress_bits_addr = _T_16 ? addr_1 : io_in_writeAddress_bits_addr; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 115:10]
  assign io_out_writeAddress_bits_len = _T_16 ? address_1_len : io_in_writeAddress_bits_len; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 115:10]
  assign io_out_writeAddress_bits_size = io_in_writeAddress_bits_size; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 115:10]
  assign io_out_writeAddress_bits_burst = io_in_writeAddress_bits_burst; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 115:10]
  assign io_out_writeAddress_bits_lock = io_in_writeAddress_bits_lock; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 115:10]
  assign io_out_writeAddress_bits_cache = io_in_writeAddress_bits_cache; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 115:10]
  assign io_out_writeAddress_bits_prot = io_in_writeAddress_bits_prot; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 115:10]
  assign io_out_writeAddress_bits_qos = io_in_writeAddress_bits_qos; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 115:10]
  assign io_out_writeData_valid = writeSplitter_io_out_valid; // @[MemBoundarySplitter.scala 128:20]
  assign io_out_writeData_bits_id = writeSplitter_io_out_bits_id; // @[MemBoundarySplitter.scala 128:20]
  assign io_out_writeData_bits_data = writeSplitter_io_out_bits_data; // @[MemBoundarySplitter.scala 128:20]
  assign io_out_writeData_bits_strb = writeSplitter_io_out_bits_strb; // @[MemBoundarySplitter.scala 128:20]
  assign io_out_writeData_bits_last = writeSplitter_io_out_bits_last; // @[MemBoundarySplitter.scala 128:20]
  assign io_out_writeResponse_ready = writeResponseFilter_io_in_ready; // @[MemBoundarySplitter.scala 131:29]
  assign io_out_readAddress_valid = _T_5 ? _GEN_22 : ready_io_out_readAddress_w_valid; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 85:10]
  assign io_out_readAddress_bits_id = io_in_readAddress_bits_id; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 85:10]
  assign io_out_readAddress_bits_addr = _T_5 ? addr : io_in_readAddress_bits_addr; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 85:10]
  assign io_out_readAddress_bits_len = _T_5 ? address_len : io_in_readAddress_bits_len; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 85:10]
  assign io_out_readAddress_bits_size = io_in_readAddress_bits_size; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 85:10]
  assign io_out_readAddress_bits_burst = io_in_readAddress_bits_burst; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 85:10]
  assign io_out_readAddress_bits_lock = io_in_readAddress_bits_lock; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 85:10]
  assign io_out_readAddress_bits_cache = io_in_readAddress_bits_cache; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 85:10]
  assign io_out_readAddress_bits_prot = io_in_readAddress_bits_prot; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 85:10]
  assign io_out_readAddress_bits_qos = io_in_readAddress_bits_qos; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 85:10]
  assign io_out_readData_ready = readMerger_io_in_ready; // @[MemBoundarySplitter.scala 123:20]
  assign readDataQueue_clock = clock;
  assign readDataQueue_reset = reset;
  assign readDataQueue_io_enq_valid = _T_5 ? _GEN_33 : ready_readDataQueue_io_enq_w_valid; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 86:10]
  assign readDataQueue_io_enq_bits = io_in_readAddress_bits_len; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 86:10]
  assign readDataQueue_io_deq_ready = readMerger_io_control_ready; // @[MemBoundarySplitter.scala 122:25]
  assign writeDataQueue_clock = clock;
  assign writeDataQueue_reset = reset;
  assign writeDataQueue_io_enq_valid = _T_16 ? _GEN_96 : ready_writeDataQueue_io_enq_w_1_valid; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 116:10]
  assign writeDataQueue_io_enq_bits = _T_16 ? address_1_len : io_in_writeAddress_bits_len; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 116:10]
  assign writeDataQueue_io_deq_ready = writeSplitter_io_control_ready; // @[MemBoundarySplitter.scala 126:28]
  assign writeResponseQueue_clock = clock;
  assign writeResponseQueue_reset = reset;
  assign writeResponseQueue_io_enq_valid = _T_16 ? _GEN_99 : ready_writeResponseQueue_io_enq_w_1_valid; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 117:10]
  assign writeResponseQueue_io_enq_bits = _T_16 ? _GEN_100 : 1'h1; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 117:10]
  assign writeResponseQueue_io_deq_ready = writeResponseFilter_io_control_ready; // @[MemBoundarySplitter.scala 130:34]
  assign readMerger_clock = clock;
  assign readMerger_reset = reset;
  assign readMerger_io_control_valid = readDataQueue_io_deq_valid; // @[MemBoundarySplitter.scala 122:25]
  assign readMerger_io_control_bits = readDataQueue_io_deq_bits; // @[MemBoundarySplitter.scala 122:25]
  assign readMerger_io_in_valid = io_out_readData_valid; // @[MemBoundarySplitter.scala 123:20]
  assign readMerger_io_in_bits_data = io_out_readData_bits_data; // @[MemBoundarySplitter.scala 123:20]
  assign readMerger_io_out_ready = io_in_readData_ready; // @[MemBoundarySplitter.scala 124:18]
  assign writeSplitter_clock = clock;
  assign writeSplitter_reset = reset;
  assign writeSplitter_io_control_valid = writeDataQueue_io_deq_valid; // @[MemBoundarySplitter.scala 126:28]
  assign writeSplitter_io_control_bits = writeDataQueue_io_deq_bits; // @[MemBoundarySplitter.scala 126:28]
  assign writeSplitter_io_in_valid = io_in_writeData_valid; // @[MemBoundarySplitter.scala 127:23]
  assign writeSplitter_io_in_bits_id = io_in_writeData_bits_id; // @[MemBoundarySplitter.scala 127:23]
  assign writeSplitter_io_in_bits_data = io_in_writeData_bits_data; // @[MemBoundarySplitter.scala 127:23]
  assign writeSplitter_io_in_bits_strb = io_in_writeData_bits_strb; // @[MemBoundarySplitter.scala 127:23]
  assign writeSplitter_io_out_ready = io_out_writeData_ready; // @[MemBoundarySplitter.scala 128:20]
  assign writeResponseFilter_io_control_valid = writeResponseQueue_io_deq_valid; // @[MemBoundarySplitter.scala 130:34]
  assign writeResponseFilter_io_control_bits = writeResponseQueue_io_deq_bits; // @[MemBoundarySplitter.scala 130:34]
  assign writeResponseFilter_io_in_valid = io_out_writeResponse_valid; // @[MemBoundarySplitter.scala 131:29]
  assign writeResponseFilter_io_out_ready = io_in_writeResponse_ready; // @[MemBoundarySplitter.scala 132:23]
  assign readEnqueuer_clock = clock;
  assign readEnqueuer_reset = reset;
  assign readEnqueuer_io_in_valid = _T_5 ? _GEN_20 : io_in_readAddress_valid; // @[MemBoundarySplitter.scala 150:74 MultiEnqueue.scala 84:17]
  assign readEnqueuer_io_out_0_ready = _T_5 ? _GEN_21 : io_out_readAddress_ready; // @[MemBoundarySplitter.scala 150:74 ReadyValid.scala 19:11]
  assign readEnqueuer_io_out_1_ready = _T_5 ? _GEN_32 : ready_readDataQueue_io_enq_w_ready; // @[MemBoundarySplitter.scala 150:74 ReadyValid.scala 19:11]
  assign writeEnqueuer_clock = clock;
  assign writeEnqueuer_reset = reset;
  assign writeEnqueuer_io_in_valid = io_in_writeAddress_valid; // @[MemBoundarySplitter.scala 224:76 MultiEnqueue.scala 114:17]
  assign writeEnqueuer_io_out_0_ready = io_out_writeAddress_ready; // @[MemBoundarySplitter.scala 224:76 ReadyValid.scala 19:11]
  assign writeEnqueuer_io_out_1_ready = _T_16 ? _GEN_95 : ready_writeDataQueue_io_enq_w_1_ready; // @[MemBoundarySplitter.scala 224:76 ReadyValid.scala 19:11]
  assign writeEnqueuer_io_out_2_ready = _T_16 ? _GEN_98 : ready_writeResponseQueue_io_enq_w_1_ready; // @[MemBoundarySplitter.scala 224:76 ReadyValid.scala 19:11]
  always @(posedge clock) begin
    readAddressCounter <= _GEN_137[11:0]; // @[MemBoundarySplitter.scala 137:{35,35}]
    readLenCounter <= _GEN_138[7:0]; // @[MemBoundarySplitter.scala 140:{31,31}]
    writeAddressCounter <= _GEN_139[11:0]; // @[MemBoundarySplitter.scala 141:{36,36}]
    writeLenCounter <= _GEN_140[7:0]; // @[MemBoundarySplitter.scala 144:{32,32}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  readAddressCounter = _RAND_0[11:0];
  _RAND_1 = {1{`RANDOM}};
  readLenCounter = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  writeAddressCounter = _RAND_2[11:0];
  _RAND_3 = {1{`RANDOM}};
  writeLenCounter = _RAND_3[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_36(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_write,
  input  [20:0] io_enq_bits_address,
  input  [20:0] io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_write,
  output [20:0] io_deq_bits_address,
  output [20:0] io_deq_bits_size
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  ram_write [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_write_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_write_MPORT_en; // @[Decoupled.scala 259:95]
  reg [20:0] ram_address [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [20:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [20:0] ram_address_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 259:95]
  reg [20:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [20:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [20:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_write_io_deq_bits_MPORT_en = 1'h1;
  assign ram_write_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_write_io_deq_bits_MPORT_data = ram_write[ram_write_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_write_MPORT_data = io_enq_bits_write;
  assign ram_write_MPORT_addr = enq_ptr_value;
  assign ram_write_MPORT_mask = 1'h1;
  assign ram_write_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = enq_ptr_value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_write = ram_write_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_write_MPORT_en & ram_write_MPORT_mask) begin
      ram_write[ram_write_MPORT_addr] <= ram_write_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_write[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_1[20:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[20:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RequestSplitter(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_write,
  input  [20:0] io_in_bits_address,
  input  [20:0] io_in_bits_size,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_write,
  output [20:0] io_out_bits_address,
  output [20:0] io_out_bits_size
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] sizeCounter; // @[RequestSplitter.scala 21:33]
  reg  sizeCounterValid; // @[RequestSplitter.scala 22:33]
  reg [20:0] addressOffset; // @[RequestSplitter.scala 23:33]
  wire [20:0] address = io_in_bits_address + addressOffset; // @[RequestSplitter.scala 24:42]
  wire  _T_3 = io_in_valid & io_out_ready; // @[RequestSplitter.scala 38:21]
  wire [20:0] _sizeCounter_T_1 = sizeCounter - 21'h40; // @[RequestSplitter.scala 53:38]
  wire [20:0] _addressOffset_T_1 = addressOffset + 21'h40; // @[RequestSplitter.scala 54:42]
  wire [20:0] _sizeCounter_T_3 = io_in_bits_size - 21'h40; // @[RequestSplitter.scala 56:39]
  wire [20:0] _GEN_2 = sizeCounterValid ? _sizeCounter_T_1 : _sizeCounter_T_3; // @[RequestSplitter.scala 52:32 53:23 56:23]
  wire [20:0] _GEN_3 = sizeCounterValid ? _addressOffset_T_1 : 21'h40; // @[RequestSplitter.scala 52:32 54:25 57:25]
  wire  _GEN_4 = sizeCounterValid ? sizeCounterValid : 1'h1; // @[RequestSplitter.scala 52:32 22:33 58:28]
  wire [20:0] _GEN_10 = sizeCounterValid & sizeCounter < 21'h40 ? sizeCounter : 21'h3f; // @[RequestSplitter.scala 29:55 30:19 43:19]
  wire  _GEN_12 = sizeCounterValid & sizeCounter < 21'h40 & io_out_ready; // @[RequestSplitter.scala 29:55 37:16 50:16]
  assign io_in_ready = io_in_bits_size < 21'h40 ? io_out_ready : _GEN_12; // @[RequestSplitter.scala 26:34 27:12]
  assign io_out_valid = io_in_valid; // @[RequestSplitter.scala 26:34 27:12]
  assign io_out_bits_write = io_in_bits_write; // @[RequestSplitter.scala 26:34 27:12]
  assign io_out_bits_address = io_in_bits_size < 21'h40 ? io_in_bits_address : address; // @[RequestSplitter.scala 26:34 27:12]
  assign io_out_bits_size = io_in_bits_size < 21'h40 ? io_in_bits_size : _GEN_10; // @[RequestSplitter.scala 26:34 27:12]
  always @(posedge clock) begin
    if (reset) begin // @[RequestSplitter.scala 21:33]
      sizeCounter <= 21'h0; // @[RequestSplitter.scala 21:33]
    end else if (!(io_in_bits_size < 21'h40)) begin // @[RequestSplitter.scala 26:34]
      if (!(sizeCounterValid & sizeCounter < 21'h40)) begin // @[RequestSplitter.scala 29:55]
        if (_T_3) begin // @[RequestSplitter.scala 51:38]
          sizeCounter <= _GEN_2;
        end
      end
    end
    if (reset) begin // @[RequestSplitter.scala 22:33]
      sizeCounterValid <= 1'h0; // @[RequestSplitter.scala 22:33]
    end else if (!(io_in_bits_size < 21'h40)) begin // @[RequestSplitter.scala 26:34]
      if (sizeCounterValid & sizeCounter < 21'h40) begin // @[RequestSplitter.scala 29:55]
        if (io_in_valid & io_out_ready) begin // @[RequestSplitter.scala 38:38]
          sizeCounterValid <= 1'h0; // @[RequestSplitter.scala 39:26]
        end
      end else if (_T_3) begin // @[RequestSplitter.scala 51:38]
        sizeCounterValid <= _GEN_4;
      end
    end
    if (reset) begin // @[RequestSplitter.scala 23:33]
      addressOffset <= 21'h0; // @[RequestSplitter.scala 23:33]
    end else if (!(io_in_bits_size < 21'h40)) begin // @[RequestSplitter.scala 26:34]
      if (sizeCounterValid & sizeCounter < 21'h40) begin // @[RequestSplitter.scala 29:55]
        if (io_in_valid & io_out_ready) begin // @[RequestSplitter.scala 38:38]
          addressOffset <= 21'h0; // @[RequestSplitter.scala 40:23]
        end
      end else if (_T_3) begin // @[RequestSplitter.scala 51:38]
        addressOffset <= _GEN_3;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sizeCounter = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  sizeCounterValid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  addressOffset = _RAND_2[20:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_37(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_0,
  input  [15:0] io_enq_bits_1,
  input  [15:0] io_enq_bits_2,
  input  [15:0] io_enq_bits_3,
  input  [15:0] io_enq_bits_4,
  input  [15:0] io_enq_bits_5,
  input  [15:0] io_enq_bits_6,
  input  [15:0] io_enq_bits_7,
  input  [15:0] io_enq_bits_8,
  input  [15:0] io_enq_bits_9,
  input  [15:0] io_enq_bits_10,
  input  [15:0] io_enq_bits_11,
  input  [15:0] io_enq_bits_12,
  input  [15:0] io_enq_bits_13,
  input  [15:0] io_enq_bits_14,
  input  [15:0] io_enq_bits_15,
  input  [15:0] io_enq_bits_16,
  input  [15:0] io_enq_bits_17,
  input  [15:0] io_enq_bits_18,
  input  [15:0] io_enq_bits_19,
  input  [15:0] io_enq_bits_20,
  input  [15:0] io_enq_bits_21,
  input  [15:0] io_enq_bits_22,
  input  [15:0] io_enq_bits_23,
  input  [15:0] io_enq_bits_24,
  input  [15:0] io_enq_bits_25,
  input  [15:0] io_enq_bits_26,
  input  [15:0] io_enq_bits_27,
  input  [15:0] io_enq_bits_28,
  input  [15:0] io_enq_bits_29,
  input  [15:0] io_enq_bits_30,
  input  [15:0] io_enq_bits_31,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_0,
  output [15:0] io_deq_bits_1,
  output [15:0] io_deq_bits_2,
  output [15:0] io_deq_bits_3,
  output [15:0] io_deq_bits_4,
  output [15:0] io_deq_bits_5,
  output [15:0] io_deq_bits_6,
  output [15:0] io_deq_bits_7,
  output [15:0] io_deq_bits_8,
  output [15:0] io_deq_bits_9,
  output [15:0] io_deq_bits_10,
  output [15:0] io_deq_bits_11,
  output [15:0] io_deq_bits_12,
  output [15:0] io_deq_bits_13,
  output [15:0] io_deq_bits_14,
  output [15:0] io_deq_bits_15,
  output [15:0] io_deq_bits_16,
  output [15:0] io_deq_bits_17,
  output [15:0] io_deq_bits_18,
  output [15:0] io_deq_bits_19,
  output [15:0] io_deq_bits_20,
  output [15:0] io_deq_bits_21,
  output [15:0] io_deq_bits_22,
  output [15:0] io_deq_bits_23,
  output [15:0] io_deq_bits_24,
  output [15:0] io_deq_bits_25,
  output [15:0] io_deq_bits_26,
  output [15:0] io_deq_bits_27,
  output [15:0] io_deq_bits_28,
  output [15:0] io_deq_bits_29,
  output [15:0] io_deq_bits_30,
  output [15:0] io_deq_bits_31
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ram_0 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_1 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_2 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_3 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_4 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_5 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_6 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_7 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_8 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_8_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_8_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_8_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_8_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_8_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_8_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_8_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_9 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_9_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_9_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_9_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_9_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_9_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_9_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_9_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_10 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_10_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_10_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_10_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_10_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_10_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_10_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_10_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_11 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_11_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_11_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_11_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_11_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_11_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_11_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_11_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_12 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_12_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_12_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_12_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_12_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_12_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_12_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_12_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_13 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_13_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_13_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_13_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_13_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_13_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_13_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_13_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_14 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_14_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_14_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_14_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_14_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_14_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_14_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_14_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_15 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_15_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_15_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_15_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_15_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_15_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_15_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_15_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_16 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_16_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_16_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_16_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_16_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_16_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_16_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_16_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_17 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_17_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_17_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_17_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_17_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_17_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_17_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_17_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_18 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_18_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_18_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_18_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_18_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_18_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_18_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_18_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_19 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_19_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_19_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_19_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_19_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_19_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_19_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_19_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_20 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_20_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_20_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_20_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_20_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_20_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_20_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_20_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_21 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_21_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_21_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_21_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_21_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_21_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_21_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_21_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_22 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_22_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_22_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_22_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_22_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_22_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_22_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_22_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_23 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_23_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_23_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_23_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_23_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_23_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_23_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_23_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_24 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_24_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_24_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_24_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_24_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_24_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_24_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_24_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_25 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_25_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_25_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_25_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_25_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_25_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_25_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_25_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_26 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_26_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_26_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_26_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_26_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_26_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_26_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_26_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_27 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_27_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_27_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_27_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_27_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_27_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_27_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_27_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_28 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_28_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_28_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_28_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_28_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_28_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_28_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_28_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_29 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_29_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_29_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_29_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_29_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_29_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_29_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_29_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_30 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_30_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_30_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_30_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_30_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_30_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_30_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_30_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_31 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_31_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_31_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_31_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_31_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_31_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_31_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_31_MPORT_en; // @[Decoupled.scala 259:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_0_io_deq_bits_MPORT_data = ram_0[ram_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_0_MPORT_data = io_enq_bits_0;
  assign ram_0_MPORT_addr = enq_ptr_value;
  assign ram_0_MPORT_mask = 1'h1;
  assign ram_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_1_io_deq_bits_MPORT_data = ram_1[ram_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_1_MPORT_data = io_enq_bits_1;
  assign ram_1_MPORT_addr = enq_ptr_value;
  assign ram_1_MPORT_mask = 1'h1;
  assign ram_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_2_io_deq_bits_MPORT_data = ram_2[ram_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_2_MPORT_data = io_enq_bits_2;
  assign ram_2_MPORT_addr = enq_ptr_value;
  assign ram_2_MPORT_mask = 1'h1;
  assign ram_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_3_io_deq_bits_MPORT_data = ram_3[ram_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_3_MPORT_data = io_enq_bits_3;
  assign ram_3_MPORT_addr = enq_ptr_value;
  assign ram_3_MPORT_mask = 1'h1;
  assign ram_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_4_io_deq_bits_MPORT_data = ram_4[ram_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_4_MPORT_data = io_enq_bits_4;
  assign ram_4_MPORT_addr = enq_ptr_value;
  assign ram_4_MPORT_mask = 1'h1;
  assign ram_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_5_io_deq_bits_MPORT_data = ram_5[ram_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_5_MPORT_data = io_enq_bits_5;
  assign ram_5_MPORT_addr = enq_ptr_value;
  assign ram_5_MPORT_mask = 1'h1;
  assign ram_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_6_io_deq_bits_MPORT_data = ram_6[ram_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_6_MPORT_data = io_enq_bits_6;
  assign ram_6_MPORT_addr = enq_ptr_value;
  assign ram_6_MPORT_mask = 1'h1;
  assign ram_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_7_io_deq_bits_MPORT_data = ram_7[ram_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_7_MPORT_data = io_enq_bits_7;
  assign ram_7_MPORT_addr = enq_ptr_value;
  assign ram_7_MPORT_mask = 1'h1;
  assign ram_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_8_io_deq_bits_MPORT_en = 1'h1;
  assign ram_8_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_8_io_deq_bits_MPORT_data = ram_8[ram_8_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_8_MPORT_data = io_enq_bits_8;
  assign ram_8_MPORT_addr = enq_ptr_value;
  assign ram_8_MPORT_mask = 1'h1;
  assign ram_8_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_9_io_deq_bits_MPORT_en = 1'h1;
  assign ram_9_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_9_io_deq_bits_MPORT_data = ram_9[ram_9_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_9_MPORT_data = io_enq_bits_9;
  assign ram_9_MPORT_addr = enq_ptr_value;
  assign ram_9_MPORT_mask = 1'h1;
  assign ram_9_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_10_io_deq_bits_MPORT_en = 1'h1;
  assign ram_10_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_10_io_deq_bits_MPORT_data = ram_10[ram_10_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_10_MPORT_data = io_enq_bits_10;
  assign ram_10_MPORT_addr = enq_ptr_value;
  assign ram_10_MPORT_mask = 1'h1;
  assign ram_10_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_11_io_deq_bits_MPORT_en = 1'h1;
  assign ram_11_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_11_io_deq_bits_MPORT_data = ram_11[ram_11_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_11_MPORT_data = io_enq_bits_11;
  assign ram_11_MPORT_addr = enq_ptr_value;
  assign ram_11_MPORT_mask = 1'h1;
  assign ram_11_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_12_io_deq_bits_MPORT_en = 1'h1;
  assign ram_12_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_12_io_deq_bits_MPORT_data = ram_12[ram_12_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_12_MPORT_data = io_enq_bits_12;
  assign ram_12_MPORT_addr = enq_ptr_value;
  assign ram_12_MPORT_mask = 1'h1;
  assign ram_12_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_13_io_deq_bits_MPORT_en = 1'h1;
  assign ram_13_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_13_io_deq_bits_MPORT_data = ram_13[ram_13_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_13_MPORT_data = io_enq_bits_13;
  assign ram_13_MPORT_addr = enq_ptr_value;
  assign ram_13_MPORT_mask = 1'h1;
  assign ram_13_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_14_io_deq_bits_MPORT_en = 1'h1;
  assign ram_14_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_14_io_deq_bits_MPORT_data = ram_14[ram_14_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_14_MPORT_data = io_enq_bits_14;
  assign ram_14_MPORT_addr = enq_ptr_value;
  assign ram_14_MPORT_mask = 1'h1;
  assign ram_14_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_15_io_deq_bits_MPORT_en = 1'h1;
  assign ram_15_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_15_io_deq_bits_MPORT_data = ram_15[ram_15_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_15_MPORT_data = io_enq_bits_15;
  assign ram_15_MPORT_addr = enq_ptr_value;
  assign ram_15_MPORT_mask = 1'h1;
  assign ram_15_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_16_io_deq_bits_MPORT_en = 1'h1;
  assign ram_16_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_16_io_deq_bits_MPORT_data = ram_16[ram_16_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_16_MPORT_data = io_enq_bits_16;
  assign ram_16_MPORT_addr = enq_ptr_value;
  assign ram_16_MPORT_mask = 1'h1;
  assign ram_16_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_17_io_deq_bits_MPORT_en = 1'h1;
  assign ram_17_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_17_io_deq_bits_MPORT_data = ram_17[ram_17_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_17_MPORT_data = io_enq_bits_17;
  assign ram_17_MPORT_addr = enq_ptr_value;
  assign ram_17_MPORT_mask = 1'h1;
  assign ram_17_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_18_io_deq_bits_MPORT_en = 1'h1;
  assign ram_18_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_18_io_deq_bits_MPORT_data = ram_18[ram_18_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_18_MPORT_data = io_enq_bits_18;
  assign ram_18_MPORT_addr = enq_ptr_value;
  assign ram_18_MPORT_mask = 1'h1;
  assign ram_18_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_19_io_deq_bits_MPORT_en = 1'h1;
  assign ram_19_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_19_io_deq_bits_MPORT_data = ram_19[ram_19_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_19_MPORT_data = io_enq_bits_19;
  assign ram_19_MPORT_addr = enq_ptr_value;
  assign ram_19_MPORT_mask = 1'h1;
  assign ram_19_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_20_io_deq_bits_MPORT_en = 1'h1;
  assign ram_20_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_20_io_deq_bits_MPORT_data = ram_20[ram_20_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_20_MPORT_data = io_enq_bits_20;
  assign ram_20_MPORT_addr = enq_ptr_value;
  assign ram_20_MPORT_mask = 1'h1;
  assign ram_20_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_21_io_deq_bits_MPORT_en = 1'h1;
  assign ram_21_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_21_io_deq_bits_MPORT_data = ram_21[ram_21_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_21_MPORT_data = io_enq_bits_21;
  assign ram_21_MPORT_addr = enq_ptr_value;
  assign ram_21_MPORT_mask = 1'h1;
  assign ram_21_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_22_io_deq_bits_MPORT_en = 1'h1;
  assign ram_22_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_22_io_deq_bits_MPORT_data = ram_22[ram_22_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_22_MPORT_data = io_enq_bits_22;
  assign ram_22_MPORT_addr = enq_ptr_value;
  assign ram_22_MPORT_mask = 1'h1;
  assign ram_22_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_23_io_deq_bits_MPORT_en = 1'h1;
  assign ram_23_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_23_io_deq_bits_MPORT_data = ram_23[ram_23_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_23_MPORT_data = io_enq_bits_23;
  assign ram_23_MPORT_addr = enq_ptr_value;
  assign ram_23_MPORT_mask = 1'h1;
  assign ram_23_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_24_io_deq_bits_MPORT_en = 1'h1;
  assign ram_24_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_24_io_deq_bits_MPORT_data = ram_24[ram_24_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_24_MPORT_data = io_enq_bits_24;
  assign ram_24_MPORT_addr = enq_ptr_value;
  assign ram_24_MPORT_mask = 1'h1;
  assign ram_24_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_25_io_deq_bits_MPORT_en = 1'h1;
  assign ram_25_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_25_io_deq_bits_MPORT_data = ram_25[ram_25_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_25_MPORT_data = io_enq_bits_25;
  assign ram_25_MPORT_addr = enq_ptr_value;
  assign ram_25_MPORT_mask = 1'h1;
  assign ram_25_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_26_io_deq_bits_MPORT_en = 1'h1;
  assign ram_26_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_26_io_deq_bits_MPORT_data = ram_26[ram_26_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_26_MPORT_data = io_enq_bits_26;
  assign ram_26_MPORT_addr = enq_ptr_value;
  assign ram_26_MPORT_mask = 1'h1;
  assign ram_26_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_27_io_deq_bits_MPORT_en = 1'h1;
  assign ram_27_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_27_io_deq_bits_MPORT_data = ram_27[ram_27_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_27_MPORT_data = io_enq_bits_27;
  assign ram_27_MPORT_addr = enq_ptr_value;
  assign ram_27_MPORT_mask = 1'h1;
  assign ram_27_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_28_io_deq_bits_MPORT_en = 1'h1;
  assign ram_28_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_28_io_deq_bits_MPORT_data = ram_28[ram_28_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_28_MPORT_data = io_enq_bits_28;
  assign ram_28_MPORT_addr = enq_ptr_value;
  assign ram_28_MPORT_mask = 1'h1;
  assign ram_28_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_29_io_deq_bits_MPORT_en = 1'h1;
  assign ram_29_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_29_io_deq_bits_MPORT_data = ram_29[ram_29_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_29_MPORT_data = io_enq_bits_29;
  assign ram_29_MPORT_addr = enq_ptr_value;
  assign ram_29_MPORT_mask = 1'h1;
  assign ram_29_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_30_io_deq_bits_MPORT_en = 1'h1;
  assign ram_30_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_30_io_deq_bits_MPORT_data = ram_30[ram_30_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_30_MPORT_data = io_enq_bits_30;
  assign ram_30_MPORT_addr = enq_ptr_value;
  assign ram_30_MPORT_mask = 1'h1;
  assign ram_30_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_31_io_deq_bits_MPORT_en = 1'h1;
  assign ram_31_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_31_io_deq_bits_MPORT_data = ram_31[ram_31_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_31_MPORT_data = io_enq_bits_31;
  assign ram_31_MPORT_addr = enq_ptr_value;
  assign ram_31_MPORT_mask = 1'h1;
  assign ram_31_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_0 = ram_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_1 = ram_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_2 = ram_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_3 = ram_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_4 = ram_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_5 = ram_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_6 = ram_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_7 = ram_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_8 = ram_8_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_9 = ram_9_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_10 = ram_10_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_11 = ram_11_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_12 = ram_12_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_13 = ram_13_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_14 = ram_14_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_15 = ram_15_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_16 = ram_16_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_17 = ram_17_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_18 = ram_18_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_19 = ram_19_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_20 = ram_20_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_21 = ram_21_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_22 = ram_22_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_23 = ram_23_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_24 = ram_24_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_25 = ram_25_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_26 = ram_26_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_27 = ram_27_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_28 = ram_28_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_29 = ram_29_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_30 = ram_30_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_31 = ram_31_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_0_MPORT_en & ram_0_MPORT_mask) begin
      ram_0[ram_0_MPORT_addr] <= ram_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_1_MPORT_en & ram_1_MPORT_mask) begin
      ram_1[ram_1_MPORT_addr] <= ram_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_2_MPORT_en & ram_2_MPORT_mask) begin
      ram_2[ram_2_MPORT_addr] <= ram_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_3_MPORT_en & ram_3_MPORT_mask) begin
      ram_3[ram_3_MPORT_addr] <= ram_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_4_MPORT_en & ram_4_MPORT_mask) begin
      ram_4[ram_4_MPORT_addr] <= ram_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_5_MPORT_en & ram_5_MPORT_mask) begin
      ram_5[ram_5_MPORT_addr] <= ram_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_6_MPORT_en & ram_6_MPORT_mask) begin
      ram_6[ram_6_MPORT_addr] <= ram_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_7_MPORT_en & ram_7_MPORT_mask) begin
      ram_7[ram_7_MPORT_addr] <= ram_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_8_MPORT_en & ram_8_MPORT_mask) begin
      ram_8[ram_8_MPORT_addr] <= ram_8_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_9_MPORT_en & ram_9_MPORT_mask) begin
      ram_9[ram_9_MPORT_addr] <= ram_9_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_10_MPORT_en & ram_10_MPORT_mask) begin
      ram_10[ram_10_MPORT_addr] <= ram_10_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_11_MPORT_en & ram_11_MPORT_mask) begin
      ram_11[ram_11_MPORT_addr] <= ram_11_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_12_MPORT_en & ram_12_MPORT_mask) begin
      ram_12[ram_12_MPORT_addr] <= ram_12_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_13_MPORT_en & ram_13_MPORT_mask) begin
      ram_13[ram_13_MPORT_addr] <= ram_13_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_14_MPORT_en & ram_14_MPORT_mask) begin
      ram_14[ram_14_MPORT_addr] <= ram_14_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_15_MPORT_en & ram_15_MPORT_mask) begin
      ram_15[ram_15_MPORT_addr] <= ram_15_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_16_MPORT_en & ram_16_MPORT_mask) begin
      ram_16[ram_16_MPORT_addr] <= ram_16_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_17_MPORT_en & ram_17_MPORT_mask) begin
      ram_17[ram_17_MPORT_addr] <= ram_17_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_18_MPORT_en & ram_18_MPORT_mask) begin
      ram_18[ram_18_MPORT_addr] <= ram_18_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_19_MPORT_en & ram_19_MPORT_mask) begin
      ram_19[ram_19_MPORT_addr] <= ram_19_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_20_MPORT_en & ram_20_MPORT_mask) begin
      ram_20[ram_20_MPORT_addr] <= ram_20_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_21_MPORT_en & ram_21_MPORT_mask) begin
      ram_21[ram_21_MPORT_addr] <= ram_21_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_22_MPORT_en & ram_22_MPORT_mask) begin
      ram_22[ram_22_MPORT_addr] <= ram_22_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_23_MPORT_en & ram_23_MPORT_mask) begin
      ram_23[ram_23_MPORT_addr] <= ram_23_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_24_MPORT_en & ram_24_MPORT_mask) begin
      ram_24[ram_24_MPORT_addr] <= ram_24_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_25_MPORT_en & ram_25_MPORT_mask) begin
      ram_25[ram_25_MPORT_addr] <= ram_25_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_26_MPORT_en & ram_26_MPORT_mask) begin
      ram_26[ram_26_MPORT_addr] <= ram_26_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_27_MPORT_en & ram_27_MPORT_mask) begin
      ram_27[ram_27_MPORT_addr] <= ram_27_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_28_MPORT_en & ram_28_MPORT_mask) begin
      ram_28[ram_28_MPORT_addr] <= ram_28_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_29_MPORT_en & ram_29_MPORT_mask) begin
      ram_29[ram_29_MPORT_addr] <= ram_29_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_30_MPORT_en & ram_30_MPORT_mask) begin
      ram_30[ram_30_MPORT_addr] <= ram_30_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_31_MPORT_en & ram_31_MPORT_mask) begin
      ram_31[ram_31_MPORT_addr] <= ram_31_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_0[initvar] = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_1[initvar] = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_2[initvar] = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_3[initvar] = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_4[initvar] = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_5[initvar] = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_6[initvar] = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_7[initvar] = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_8[initvar] = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_9[initvar] = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_10[initvar] = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_11[initvar] = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_12[initvar] = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_13[initvar] = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_14[initvar] = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_15[initvar] = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_16[initvar] = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_17[initvar] = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_18[initvar] = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_19[initvar] = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_20[initvar] = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_21[initvar] = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_22[initvar] = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_23[initvar] = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_24[initvar] = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_25[initvar] = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_26[initvar] = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_27[initvar] = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_28[initvar] = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_29[initvar] = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_30[initvar] = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_31[initvar] = _RAND_31[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  enq_ptr_value = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  deq_ptr_value = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  maybe_full = _RAND_34[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_38(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits_data,
  input          io_enq_bits_last,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits_data,
  output         io_deq_bits_last
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [127:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [127:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_last [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 259:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = enq_ptr_value;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[127:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = _RAND_1[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_39(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_deq_ready,
  output  io_deq_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enq_ptr_value = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  deq_ptr_value = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module VectorSerializer(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [15:0]  io_in_bits_0,
  input  [15:0]  io_in_bits_1,
  input  [15:0]  io_in_bits_2,
  input  [15:0]  io_in_bits_3,
  input  [15:0]  io_in_bits_4,
  input  [15:0]  io_in_bits_5,
  input  [15:0]  io_in_bits_6,
  input  [15:0]  io_in_bits_7,
  input  [15:0]  io_in_bits_8,
  input  [15:0]  io_in_bits_9,
  input  [15:0]  io_in_bits_10,
  input  [15:0]  io_in_bits_11,
  input  [15:0]  io_in_bits_12,
  input  [15:0]  io_in_bits_13,
  input  [15:0]  io_in_bits_14,
  input  [15:0]  io_in_bits_15,
  input  [15:0]  io_in_bits_16,
  input  [15:0]  io_in_bits_17,
  input  [15:0]  io_in_bits_18,
  input  [15:0]  io_in_bits_19,
  input  [15:0]  io_in_bits_20,
  input  [15:0]  io_in_bits_21,
  input  [15:0]  io_in_bits_22,
  input  [15:0]  io_in_bits_23,
  input  [15:0]  io_in_bits_24,
  input  [15:0]  io_in_bits_25,
  input  [15:0]  io_in_bits_26,
  input  [15:0]  io_in_bits_27,
  input  [15:0]  io_in_bits_28,
  input  [15:0]  io_in_bits_29,
  input  [15:0]  io_in_bits_30,
  input  [15:0]  io_in_bits_31,
  input          io_out_ready,
  output         io_out_valid,
  output [127:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] bits_0; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_1; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_2; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_3; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_4; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_5; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_6; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_7; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_8; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_9; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_10; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_11; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_12; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_13; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_14; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_15; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_16; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_17; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_18; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_19; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_20; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_21; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_22; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_23; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_24; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_25; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_26; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_27; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_28; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_29; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_30; // @[VectorSerializer.scala 37:22]
  reg [15:0] bits_31; // @[VectorSerializer.scala 37:22]
  reg  valid; // @[VectorSerializer.scala 38:22]
  wire  _T = valid & io_out_ready; // @[VectorSerializer.scala 40:48]
  reg [1:0] ctr; // @[Counter.scala 62:40]
  wire  wrap_wrap = ctr == 2'h3; // @[Counter.scala 74:24]
  wire [1:0] _wrap_value_T_1 = ctr + 2'h1; // @[Counter.scala 78:24]
  wire  wrap = _T & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire [5:0] _out_T = ctr * 4'h8; // @[VectorSerializer.scala 46:18]
  wire [6:0] _out_T_1 = {{1'd0}, _out_T}; // @[VectorSerializer.scala 46:40]
  wire [15:0] _GEN_3 = 5'h1 == _out_T_1[4:0] ? $signed(bits_1) : $signed(bits_0); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_4 = 5'h2 == _out_T_1[4:0] ? $signed(bits_2) : $signed(_GEN_3); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_5 = 5'h3 == _out_T_1[4:0] ? $signed(bits_3) : $signed(_GEN_4); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_6 = 5'h4 == _out_T_1[4:0] ? $signed(bits_4) : $signed(_GEN_5); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_7 = 5'h5 == _out_T_1[4:0] ? $signed(bits_5) : $signed(_GEN_6); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_8 = 5'h6 == _out_T_1[4:0] ? $signed(bits_6) : $signed(_GEN_7); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_9 = 5'h7 == _out_T_1[4:0] ? $signed(bits_7) : $signed(_GEN_8); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_10 = 5'h8 == _out_T_1[4:0] ? $signed(bits_8) : $signed(_GEN_9); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_11 = 5'h9 == _out_T_1[4:0] ? $signed(bits_9) : $signed(_GEN_10); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_12 = 5'ha == _out_T_1[4:0] ? $signed(bits_10) : $signed(_GEN_11); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_13 = 5'hb == _out_T_1[4:0] ? $signed(bits_11) : $signed(_GEN_12); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_14 = 5'hc == _out_T_1[4:0] ? $signed(bits_12) : $signed(_GEN_13); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_15 = 5'hd == _out_T_1[4:0] ? $signed(bits_13) : $signed(_GEN_14); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_16 = 5'he == _out_T_1[4:0] ? $signed(bits_14) : $signed(_GEN_15); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_17 = 5'hf == _out_T_1[4:0] ? $signed(bits_15) : $signed(_GEN_16); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_18 = 5'h10 == _out_T_1[4:0] ? $signed(bits_16) : $signed(_GEN_17); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_19 = 5'h11 == _out_T_1[4:0] ? $signed(bits_17) : $signed(_GEN_18); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_20 = 5'h12 == _out_T_1[4:0] ? $signed(bits_18) : $signed(_GEN_19); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_21 = 5'h13 == _out_T_1[4:0] ? $signed(bits_19) : $signed(_GEN_20); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_22 = 5'h14 == _out_T_1[4:0] ? $signed(bits_20) : $signed(_GEN_21); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_23 = 5'h15 == _out_T_1[4:0] ? $signed(bits_21) : $signed(_GEN_22); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_24 = 5'h16 == _out_T_1[4:0] ? $signed(bits_22) : $signed(_GEN_23); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_25 = 5'h17 == _out_T_1[4:0] ? $signed(bits_23) : $signed(_GEN_24); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_26 = 5'h18 == _out_T_1[4:0] ? $signed(bits_24) : $signed(_GEN_25); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_27 = 5'h19 == _out_T_1[4:0] ? $signed(bits_25) : $signed(_GEN_26); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_28 = 5'h1a == _out_T_1[4:0] ? $signed(bits_26) : $signed(_GEN_27); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_29 = 5'h1b == _out_T_1[4:0] ? $signed(bits_27) : $signed(_GEN_28); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_30 = 5'h1c == _out_T_1[4:0] ? $signed(bits_28) : $signed(_GEN_29); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_31 = 5'h1d == _out_T_1[4:0] ? $signed(bits_29) : $signed(_GEN_30); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_32 = 5'h1e == _out_T_1[4:0] ? $signed(bits_30) : $signed(_GEN_31); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] out_0 = 5'h1f == _out_T_1[4:0] ? $signed(bits_31) : $signed(_GEN_32); // @[VectorSerializer.scala 46:47]
  wire [5:0] _out_T_7 = _out_T + 6'h1; // @[VectorSerializer.scala 46:40]
  wire [15:0] _GEN_35 = 5'h1 == _out_T_7[4:0] ? $signed(bits_1) : $signed(bits_0); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_36 = 5'h2 == _out_T_7[4:0] ? $signed(bits_2) : $signed(_GEN_35); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_37 = 5'h3 == _out_T_7[4:0] ? $signed(bits_3) : $signed(_GEN_36); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_38 = 5'h4 == _out_T_7[4:0] ? $signed(bits_4) : $signed(_GEN_37); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_39 = 5'h5 == _out_T_7[4:0] ? $signed(bits_5) : $signed(_GEN_38); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_40 = 5'h6 == _out_T_7[4:0] ? $signed(bits_6) : $signed(_GEN_39); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_41 = 5'h7 == _out_T_7[4:0] ? $signed(bits_7) : $signed(_GEN_40); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_42 = 5'h8 == _out_T_7[4:0] ? $signed(bits_8) : $signed(_GEN_41); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_43 = 5'h9 == _out_T_7[4:0] ? $signed(bits_9) : $signed(_GEN_42); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_44 = 5'ha == _out_T_7[4:0] ? $signed(bits_10) : $signed(_GEN_43); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_45 = 5'hb == _out_T_7[4:0] ? $signed(bits_11) : $signed(_GEN_44); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_46 = 5'hc == _out_T_7[4:0] ? $signed(bits_12) : $signed(_GEN_45); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_47 = 5'hd == _out_T_7[4:0] ? $signed(bits_13) : $signed(_GEN_46); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_48 = 5'he == _out_T_7[4:0] ? $signed(bits_14) : $signed(_GEN_47); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_49 = 5'hf == _out_T_7[4:0] ? $signed(bits_15) : $signed(_GEN_48); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_50 = 5'h10 == _out_T_7[4:0] ? $signed(bits_16) : $signed(_GEN_49); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_51 = 5'h11 == _out_T_7[4:0] ? $signed(bits_17) : $signed(_GEN_50); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_52 = 5'h12 == _out_T_7[4:0] ? $signed(bits_18) : $signed(_GEN_51); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_53 = 5'h13 == _out_T_7[4:0] ? $signed(bits_19) : $signed(_GEN_52); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_54 = 5'h14 == _out_T_7[4:0] ? $signed(bits_20) : $signed(_GEN_53); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_55 = 5'h15 == _out_T_7[4:0] ? $signed(bits_21) : $signed(_GEN_54); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_56 = 5'h16 == _out_T_7[4:0] ? $signed(bits_22) : $signed(_GEN_55); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_57 = 5'h17 == _out_T_7[4:0] ? $signed(bits_23) : $signed(_GEN_56); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_58 = 5'h18 == _out_T_7[4:0] ? $signed(bits_24) : $signed(_GEN_57); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_59 = 5'h19 == _out_T_7[4:0] ? $signed(bits_25) : $signed(_GEN_58); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_60 = 5'h1a == _out_T_7[4:0] ? $signed(bits_26) : $signed(_GEN_59); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_61 = 5'h1b == _out_T_7[4:0] ? $signed(bits_27) : $signed(_GEN_60); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_62 = 5'h1c == _out_T_7[4:0] ? $signed(bits_28) : $signed(_GEN_61); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_63 = 5'h1d == _out_T_7[4:0] ? $signed(bits_29) : $signed(_GEN_62); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_64 = 5'h1e == _out_T_7[4:0] ? $signed(bits_30) : $signed(_GEN_63); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] out_1 = 5'h1f == _out_T_7[4:0] ? $signed(bits_31) : $signed(_GEN_64); // @[VectorSerializer.scala 46:47]
  wire [5:0] _out_T_12 = _out_T + 6'h2; // @[VectorSerializer.scala 46:40]
  wire [15:0] _GEN_67 = 5'h1 == _out_T_12[4:0] ? $signed(bits_1) : $signed(bits_0); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_68 = 5'h2 == _out_T_12[4:0] ? $signed(bits_2) : $signed(_GEN_67); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_69 = 5'h3 == _out_T_12[4:0] ? $signed(bits_3) : $signed(_GEN_68); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_70 = 5'h4 == _out_T_12[4:0] ? $signed(bits_4) : $signed(_GEN_69); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_71 = 5'h5 == _out_T_12[4:0] ? $signed(bits_5) : $signed(_GEN_70); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_72 = 5'h6 == _out_T_12[4:0] ? $signed(bits_6) : $signed(_GEN_71); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_73 = 5'h7 == _out_T_12[4:0] ? $signed(bits_7) : $signed(_GEN_72); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_74 = 5'h8 == _out_T_12[4:0] ? $signed(bits_8) : $signed(_GEN_73); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_75 = 5'h9 == _out_T_12[4:0] ? $signed(bits_9) : $signed(_GEN_74); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_76 = 5'ha == _out_T_12[4:0] ? $signed(bits_10) : $signed(_GEN_75); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_77 = 5'hb == _out_T_12[4:0] ? $signed(bits_11) : $signed(_GEN_76); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_78 = 5'hc == _out_T_12[4:0] ? $signed(bits_12) : $signed(_GEN_77); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_79 = 5'hd == _out_T_12[4:0] ? $signed(bits_13) : $signed(_GEN_78); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_80 = 5'he == _out_T_12[4:0] ? $signed(bits_14) : $signed(_GEN_79); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_81 = 5'hf == _out_T_12[4:0] ? $signed(bits_15) : $signed(_GEN_80); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_82 = 5'h10 == _out_T_12[4:0] ? $signed(bits_16) : $signed(_GEN_81); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_83 = 5'h11 == _out_T_12[4:0] ? $signed(bits_17) : $signed(_GEN_82); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_84 = 5'h12 == _out_T_12[4:0] ? $signed(bits_18) : $signed(_GEN_83); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_85 = 5'h13 == _out_T_12[4:0] ? $signed(bits_19) : $signed(_GEN_84); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_86 = 5'h14 == _out_T_12[4:0] ? $signed(bits_20) : $signed(_GEN_85); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_87 = 5'h15 == _out_T_12[4:0] ? $signed(bits_21) : $signed(_GEN_86); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_88 = 5'h16 == _out_T_12[4:0] ? $signed(bits_22) : $signed(_GEN_87); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_89 = 5'h17 == _out_T_12[4:0] ? $signed(bits_23) : $signed(_GEN_88); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_90 = 5'h18 == _out_T_12[4:0] ? $signed(bits_24) : $signed(_GEN_89); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_91 = 5'h19 == _out_T_12[4:0] ? $signed(bits_25) : $signed(_GEN_90); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_92 = 5'h1a == _out_T_12[4:0] ? $signed(bits_26) : $signed(_GEN_91); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_93 = 5'h1b == _out_T_12[4:0] ? $signed(bits_27) : $signed(_GEN_92); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_94 = 5'h1c == _out_T_12[4:0] ? $signed(bits_28) : $signed(_GEN_93); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_95 = 5'h1d == _out_T_12[4:0] ? $signed(bits_29) : $signed(_GEN_94); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_96 = 5'h1e == _out_T_12[4:0] ? $signed(bits_30) : $signed(_GEN_95); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] out_2 = 5'h1f == _out_T_12[4:0] ? $signed(bits_31) : $signed(_GEN_96); // @[VectorSerializer.scala 46:47]
  wire [5:0] _out_T_17 = _out_T + 6'h3; // @[VectorSerializer.scala 46:40]
  wire [15:0] _GEN_99 = 5'h1 == _out_T_17[4:0] ? $signed(bits_1) : $signed(bits_0); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_100 = 5'h2 == _out_T_17[4:0] ? $signed(bits_2) : $signed(_GEN_99); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_101 = 5'h3 == _out_T_17[4:0] ? $signed(bits_3) : $signed(_GEN_100); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_102 = 5'h4 == _out_T_17[4:0] ? $signed(bits_4) : $signed(_GEN_101); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_103 = 5'h5 == _out_T_17[4:0] ? $signed(bits_5) : $signed(_GEN_102); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_104 = 5'h6 == _out_T_17[4:0] ? $signed(bits_6) : $signed(_GEN_103); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_105 = 5'h7 == _out_T_17[4:0] ? $signed(bits_7) : $signed(_GEN_104); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_106 = 5'h8 == _out_T_17[4:0] ? $signed(bits_8) : $signed(_GEN_105); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_107 = 5'h9 == _out_T_17[4:0] ? $signed(bits_9) : $signed(_GEN_106); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_108 = 5'ha == _out_T_17[4:0] ? $signed(bits_10) : $signed(_GEN_107); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_109 = 5'hb == _out_T_17[4:0] ? $signed(bits_11) : $signed(_GEN_108); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_110 = 5'hc == _out_T_17[4:0] ? $signed(bits_12) : $signed(_GEN_109); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_111 = 5'hd == _out_T_17[4:0] ? $signed(bits_13) : $signed(_GEN_110); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_112 = 5'he == _out_T_17[4:0] ? $signed(bits_14) : $signed(_GEN_111); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_113 = 5'hf == _out_T_17[4:0] ? $signed(bits_15) : $signed(_GEN_112); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_114 = 5'h10 == _out_T_17[4:0] ? $signed(bits_16) : $signed(_GEN_113); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_115 = 5'h11 == _out_T_17[4:0] ? $signed(bits_17) : $signed(_GEN_114); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_116 = 5'h12 == _out_T_17[4:0] ? $signed(bits_18) : $signed(_GEN_115); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_117 = 5'h13 == _out_T_17[4:0] ? $signed(bits_19) : $signed(_GEN_116); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_118 = 5'h14 == _out_T_17[4:0] ? $signed(bits_20) : $signed(_GEN_117); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_119 = 5'h15 == _out_T_17[4:0] ? $signed(bits_21) : $signed(_GEN_118); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_120 = 5'h16 == _out_T_17[4:0] ? $signed(bits_22) : $signed(_GEN_119); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_121 = 5'h17 == _out_T_17[4:0] ? $signed(bits_23) : $signed(_GEN_120); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_122 = 5'h18 == _out_T_17[4:0] ? $signed(bits_24) : $signed(_GEN_121); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_123 = 5'h19 == _out_T_17[4:0] ? $signed(bits_25) : $signed(_GEN_122); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_124 = 5'h1a == _out_T_17[4:0] ? $signed(bits_26) : $signed(_GEN_123); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_125 = 5'h1b == _out_T_17[4:0] ? $signed(bits_27) : $signed(_GEN_124); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_126 = 5'h1c == _out_T_17[4:0] ? $signed(bits_28) : $signed(_GEN_125); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_127 = 5'h1d == _out_T_17[4:0] ? $signed(bits_29) : $signed(_GEN_126); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_128 = 5'h1e == _out_T_17[4:0] ? $signed(bits_30) : $signed(_GEN_127); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] out_3 = 5'h1f == _out_T_17[4:0] ? $signed(bits_31) : $signed(_GEN_128); // @[VectorSerializer.scala 46:47]
  wire [5:0] _out_T_22 = _out_T + 6'h4; // @[VectorSerializer.scala 46:40]
  wire [15:0] _GEN_131 = 5'h1 == _out_T_22[4:0] ? $signed(bits_1) : $signed(bits_0); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_132 = 5'h2 == _out_T_22[4:0] ? $signed(bits_2) : $signed(_GEN_131); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_133 = 5'h3 == _out_T_22[4:0] ? $signed(bits_3) : $signed(_GEN_132); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_134 = 5'h4 == _out_T_22[4:0] ? $signed(bits_4) : $signed(_GEN_133); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_135 = 5'h5 == _out_T_22[4:0] ? $signed(bits_5) : $signed(_GEN_134); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_136 = 5'h6 == _out_T_22[4:0] ? $signed(bits_6) : $signed(_GEN_135); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_137 = 5'h7 == _out_T_22[4:0] ? $signed(bits_7) : $signed(_GEN_136); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_138 = 5'h8 == _out_T_22[4:0] ? $signed(bits_8) : $signed(_GEN_137); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_139 = 5'h9 == _out_T_22[4:0] ? $signed(bits_9) : $signed(_GEN_138); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_140 = 5'ha == _out_T_22[4:0] ? $signed(bits_10) : $signed(_GEN_139); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_141 = 5'hb == _out_T_22[4:0] ? $signed(bits_11) : $signed(_GEN_140); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_142 = 5'hc == _out_T_22[4:0] ? $signed(bits_12) : $signed(_GEN_141); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_143 = 5'hd == _out_T_22[4:0] ? $signed(bits_13) : $signed(_GEN_142); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_144 = 5'he == _out_T_22[4:0] ? $signed(bits_14) : $signed(_GEN_143); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_145 = 5'hf == _out_T_22[4:0] ? $signed(bits_15) : $signed(_GEN_144); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_146 = 5'h10 == _out_T_22[4:0] ? $signed(bits_16) : $signed(_GEN_145); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_147 = 5'h11 == _out_T_22[4:0] ? $signed(bits_17) : $signed(_GEN_146); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_148 = 5'h12 == _out_T_22[4:0] ? $signed(bits_18) : $signed(_GEN_147); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_149 = 5'h13 == _out_T_22[4:0] ? $signed(bits_19) : $signed(_GEN_148); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_150 = 5'h14 == _out_T_22[4:0] ? $signed(bits_20) : $signed(_GEN_149); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_151 = 5'h15 == _out_T_22[4:0] ? $signed(bits_21) : $signed(_GEN_150); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_152 = 5'h16 == _out_T_22[4:0] ? $signed(bits_22) : $signed(_GEN_151); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_153 = 5'h17 == _out_T_22[4:0] ? $signed(bits_23) : $signed(_GEN_152); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_154 = 5'h18 == _out_T_22[4:0] ? $signed(bits_24) : $signed(_GEN_153); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_155 = 5'h19 == _out_T_22[4:0] ? $signed(bits_25) : $signed(_GEN_154); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_156 = 5'h1a == _out_T_22[4:0] ? $signed(bits_26) : $signed(_GEN_155); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_157 = 5'h1b == _out_T_22[4:0] ? $signed(bits_27) : $signed(_GEN_156); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_158 = 5'h1c == _out_T_22[4:0] ? $signed(bits_28) : $signed(_GEN_157); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_159 = 5'h1d == _out_T_22[4:0] ? $signed(bits_29) : $signed(_GEN_158); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_160 = 5'h1e == _out_T_22[4:0] ? $signed(bits_30) : $signed(_GEN_159); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] out_4 = 5'h1f == _out_T_22[4:0] ? $signed(bits_31) : $signed(_GEN_160); // @[VectorSerializer.scala 46:47]
  wire [5:0] _out_T_27 = _out_T + 6'h5; // @[VectorSerializer.scala 46:40]
  wire [15:0] _GEN_163 = 5'h1 == _out_T_27[4:0] ? $signed(bits_1) : $signed(bits_0); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_164 = 5'h2 == _out_T_27[4:0] ? $signed(bits_2) : $signed(_GEN_163); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_165 = 5'h3 == _out_T_27[4:0] ? $signed(bits_3) : $signed(_GEN_164); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_166 = 5'h4 == _out_T_27[4:0] ? $signed(bits_4) : $signed(_GEN_165); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_167 = 5'h5 == _out_T_27[4:0] ? $signed(bits_5) : $signed(_GEN_166); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_168 = 5'h6 == _out_T_27[4:0] ? $signed(bits_6) : $signed(_GEN_167); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_169 = 5'h7 == _out_T_27[4:0] ? $signed(bits_7) : $signed(_GEN_168); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_170 = 5'h8 == _out_T_27[4:0] ? $signed(bits_8) : $signed(_GEN_169); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_171 = 5'h9 == _out_T_27[4:0] ? $signed(bits_9) : $signed(_GEN_170); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_172 = 5'ha == _out_T_27[4:0] ? $signed(bits_10) : $signed(_GEN_171); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_173 = 5'hb == _out_T_27[4:0] ? $signed(bits_11) : $signed(_GEN_172); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_174 = 5'hc == _out_T_27[4:0] ? $signed(bits_12) : $signed(_GEN_173); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_175 = 5'hd == _out_T_27[4:0] ? $signed(bits_13) : $signed(_GEN_174); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_176 = 5'he == _out_T_27[4:0] ? $signed(bits_14) : $signed(_GEN_175); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_177 = 5'hf == _out_T_27[4:0] ? $signed(bits_15) : $signed(_GEN_176); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_178 = 5'h10 == _out_T_27[4:0] ? $signed(bits_16) : $signed(_GEN_177); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_179 = 5'h11 == _out_T_27[4:0] ? $signed(bits_17) : $signed(_GEN_178); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_180 = 5'h12 == _out_T_27[4:0] ? $signed(bits_18) : $signed(_GEN_179); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_181 = 5'h13 == _out_T_27[4:0] ? $signed(bits_19) : $signed(_GEN_180); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_182 = 5'h14 == _out_T_27[4:0] ? $signed(bits_20) : $signed(_GEN_181); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_183 = 5'h15 == _out_T_27[4:0] ? $signed(bits_21) : $signed(_GEN_182); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_184 = 5'h16 == _out_T_27[4:0] ? $signed(bits_22) : $signed(_GEN_183); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_185 = 5'h17 == _out_T_27[4:0] ? $signed(bits_23) : $signed(_GEN_184); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_186 = 5'h18 == _out_T_27[4:0] ? $signed(bits_24) : $signed(_GEN_185); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_187 = 5'h19 == _out_T_27[4:0] ? $signed(bits_25) : $signed(_GEN_186); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_188 = 5'h1a == _out_T_27[4:0] ? $signed(bits_26) : $signed(_GEN_187); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_189 = 5'h1b == _out_T_27[4:0] ? $signed(bits_27) : $signed(_GEN_188); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_190 = 5'h1c == _out_T_27[4:0] ? $signed(bits_28) : $signed(_GEN_189); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_191 = 5'h1d == _out_T_27[4:0] ? $signed(bits_29) : $signed(_GEN_190); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_192 = 5'h1e == _out_T_27[4:0] ? $signed(bits_30) : $signed(_GEN_191); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] out_5 = 5'h1f == _out_T_27[4:0] ? $signed(bits_31) : $signed(_GEN_192); // @[VectorSerializer.scala 46:47]
  wire [5:0] _out_T_32 = _out_T + 6'h6; // @[VectorSerializer.scala 46:40]
  wire [15:0] _GEN_195 = 5'h1 == _out_T_32[4:0] ? $signed(bits_1) : $signed(bits_0); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_196 = 5'h2 == _out_T_32[4:0] ? $signed(bits_2) : $signed(_GEN_195); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_197 = 5'h3 == _out_T_32[4:0] ? $signed(bits_3) : $signed(_GEN_196); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_198 = 5'h4 == _out_T_32[4:0] ? $signed(bits_4) : $signed(_GEN_197); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_199 = 5'h5 == _out_T_32[4:0] ? $signed(bits_5) : $signed(_GEN_198); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_200 = 5'h6 == _out_T_32[4:0] ? $signed(bits_6) : $signed(_GEN_199); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_201 = 5'h7 == _out_T_32[4:0] ? $signed(bits_7) : $signed(_GEN_200); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_202 = 5'h8 == _out_T_32[4:0] ? $signed(bits_8) : $signed(_GEN_201); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_203 = 5'h9 == _out_T_32[4:0] ? $signed(bits_9) : $signed(_GEN_202); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_204 = 5'ha == _out_T_32[4:0] ? $signed(bits_10) : $signed(_GEN_203); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_205 = 5'hb == _out_T_32[4:0] ? $signed(bits_11) : $signed(_GEN_204); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_206 = 5'hc == _out_T_32[4:0] ? $signed(bits_12) : $signed(_GEN_205); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_207 = 5'hd == _out_T_32[4:0] ? $signed(bits_13) : $signed(_GEN_206); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_208 = 5'he == _out_T_32[4:0] ? $signed(bits_14) : $signed(_GEN_207); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_209 = 5'hf == _out_T_32[4:0] ? $signed(bits_15) : $signed(_GEN_208); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_210 = 5'h10 == _out_T_32[4:0] ? $signed(bits_16) : $signed(_GEN_209); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_211 = 5'h11 == _out_T_32[4:0] ? $signed(bits_17) : $signed(_GEN_210); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_212 = 5'h12 == _out_T_32[4:0] ? $signed(bits_18) : $signed(_GEN_211); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_213 = 5'h13 == _out_T_32[4:0] ? $signed(bits_19) : $signed(_GEN_212); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_214 = 5'h14 == _out_T_32[4:0] ? $signed(bits_20) : $signed(_GEN_213); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_215 = 5'h15 == _out_T_32[4:0] ? $signed(bits_21) : $signed(_GEN_214); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_216 = 5'h16 == _out_T_32[4:0] ? $signed(bits_22) : $signed(_GEN_215); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_217 = 5'h17 == _out_T_32[4:0] ? $signed(bits_23) : $signed(_GEN_216); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_218 = 5'h18 == _out_T_32[4:0] ? $signed(bits_24) : $signed(_GEN_217); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_219 = 5'h19 == _out_T_32[4:0] ? $signed(bits_25) : $signed(_GEN_218); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_220 = 5'h1a == _out_T_32[4:0] ? $signed(bits_26) : $signed(_GEN_219); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_221 = 5'h1b == _out_T_32[4:0] ? $signed(bits_27) : $signed(_GEN_220); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_222 = 5'h1c == _out_T_32[4:0] ? $signed(bits_28) : $signed(_GEN_221); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_223 = 5'h1d == _out_T_32[4:0] ? $signed(bits_29) : $signed(_GEN_222); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_224 = 5'h1e == _out_T_32[4:0] ? $signed(bits_30) : $signed(_GEN_223); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] out_6 = 5'h1f == _out_T_32[4:0] ? $signed(bits_31) : $signed(_GEN_224); // @[VectorSerializer.scala 46:47]
  wire [5:0] _out_T_37 = _out_T + 6'h7; // @[VectorSerializer.scala 46:40]
  wire [15:0] _GEN_227 = 5'h1 == _out_T_37[4:0] ? $signed(bits_1) : $signed(bits_0); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_228 = 5'h2 == _out_T_37[4:0] ? $signed(bits_2) : $signed(_GEN_227); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_229 = 5'h3 == _out_T_37[4:0] ? $signed(bits_3) : $signed(_GEN_228); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_230 = 5'h4 == _out_T_37[4:0] ? $signed(bits_4) : $signed(_GEN_229); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_231 = 5'h5 == _out_T_37[4:0] ? $signed(bits_5) : $signed(_GEN_230); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_232 = 5'h6 == _out_T_37[4:0] ? $signed(bits_6) : $signed(_GEN_231); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_233 = 5'h7 == _out_T_37[4:0] ? $signed(bits_7) : $signed(_GEN_232); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_234 = 5'h8 == _out_T_37[4:0] ? $signed(bits_8) : $signed(_GEN_233); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_235 = 5'h9 == _out_T_37[4:0] ? $signed(bits_9) : $signed(_GEN_234); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_236 = 5'ha == _out_T_37[4:0] ? $signed(bits_10) : $signed(_GEN_235); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_237 = 5'hb == _out_T_37[4:0] ? $signed(bits_11) : $signed(_GEN_236); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_238 = 5'hc == _out_T_37[4:0] ? $signed(bits_12) : $signed(_GEN_237); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_239 = 5'hd == _out_T_37[4:0] ? $signed(bits_13) : $signed(_GEN_238); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_240 = 5'he == _out_T_37[4:0] ? $signed(bits_14) : $signed(_GEN_239); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_241 = 5'hf == _out_T_37[4:0] ? $signed(bits_15) : $signed(_GEN_240); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_242 = 5'h10 == _out_T_37[4:0] ? $signed(bits_16) : $signed(_GEN_241); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_243 = 5'h11 == _out_T_37[4:0] ? $signed(bits_17) : $signed(_GEN_242); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_244 = 5'h12 == _out_T_37[4:0] ? $signed(bits_18) : $signed(_GEN_243); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_245 = 5'h13 == _out_T_37[4:0] ? $signed(bits_19) : $signed(_GEN_244); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_246 = 5'h14 == _out_T_37[4:0] ? $signed(bits_20) : $signed(_GEN_245); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_247 = 5'h15 == _out_T_37[4:0] ? $signed(bits_21) : $signed(_GEN_246); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_248 = 5'h16 == _out_T_37[4:0] ? $signed(bits_22) : $signed(_GEN_247); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_249 = 5'h17 == _out_T_37[4:0] ? $signed(bits_23) : $signed(_GEN_248); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_250 = 5'h18 == _out_T_37[4:0] ? $signed(bits_24) : $signed(_GEN_249); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_251 = 5'h19 == _out_T_37[4:0] ? $signed(bits_25) : $signed(_GEN_250); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_252 = 5'h1a == _out_T_37[4:0] ? $signed(bits_26) : $signed(_GEN_251); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_253 = 5'h1b == _out_T_37[4:0] ? $signed(bits_27) : $signed(_GEN_252); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_254 = 5'h1c == _out_T_37[4:0] ? $signed(bits_28) : $signed(_GEN_253); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_255 = 5'h1d == _out_T_37[4:0] ? $signed(bits_29) : $signed(_GEN_254); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] _GEN_256 = 5'h1e == _out_T_37[4:0] ? $signed(bits_30) : $signed(_GEN_255); // @[VectorSerializer.scala 46:{47,47}]
  wire [15:0] out_7 = 5'h1f == _out_T_37[4:0] ? $signed(bits_31) : $signed(_GEN_256); // @[VectorSerializer.scala 46:47]
  wire [63:0] io_out_bits_lo = {out_3,out_2,out_1,out_0}; // @[Cat.scala 31:58]
  wire [63:0] io_out_bits_hi = {out_7,out_6,out_5,out_4}; // @[Cat.scala 31:58]
  wire [127:0] lo_lo = {io_in_bits_7,io_in_bits_6,io_in_bits_5,io_in_bits_4,io_in_bits_3,io_in_bits_2,io_in_bits_1,
    io_in_bits_0}; // @[VectorSerializer.scala 56:34]
  wire [255:0] lo = {io_in_bits_15,io_in_bits_14,io_in_bits_13,io_in_bits_12,io_in_bits_11,io_in_bits_10,io_in_bits_9,
    io_in_bits_8,lo_lo}; // @[VectorSerializer.scala 56:34]
  wire [127:0] hi_lo = {io_in_bits_23,io_in_bits_22,io_in_bits_21,io_in_bits_20,io_in_bits_19,io_in_bits_18,
    io_in_bits_17,io_in_bits_16}; // @[VectorSerializer.scala 56:34]
  wire [511:0] _T_33 = {io_in_bits_31,io_in_bits_30,io_in_bits_29,io_in_bits_28,io_in_bits_27,io_in_bits_26,
    io_in_bits_25,io_in_bits_24,hi_lo,lo}; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_35 = _T_33[15:0]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_37 = _T_33[31:16]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_39 = _T_33[47:32]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_41 = _T_33[63:48]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_43 = _T_33[79:64]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_45 = _T_33[95:80]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_47 = _T_33[111:96]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_49 = _T_33[127:112]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_51 = _T_33[143:128]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_53 = _T_33[159:144]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_55 = _T_33[175:160]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_57 = _T_33[191:176]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_59 = _T_33[207:192]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_61 = _T_33[223:208]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_63 = _T_33[239:224]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_65 = _T_33[255:240]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_67 = _T_33[271:256]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_69 = _T_33[287:272]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_71 = _T_33[303:288]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_73 = _T_33[319:304]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_75 = _T_33[335:320]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_77 = _T_33[351:336]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_79 = _T_33[367:352]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_81 = _T_33[383:368]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_83 = _T_33[399:384]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_85 = _T_33[415:400]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_87 = _T_33[431:416]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_89 = _T_33[447:432]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_91 = _T_33[463:448]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_93 = _T_33[479:464]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_95 = _T_33[495:480]; // @[VectorSerializer.scala 56:34]
  wire [15:0] _T_97 = _T_33[511:496]; // @[VectorSerializer.scala 56:34]
  assign io_in_ready = ~valid | wrap; // @[VectorSerializer.scala 52:25]
  assign io_out_valid = valid; // @[VectorSerializer.scala 50:16]
  assign io_out_bits = {io_out_bits_hi,io_out_bits_lo}; // @[Cat.scala 31:58]
  always @(posedge clock) begin
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_0 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_0 <= _T_35; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_1 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_1 <= _T_37; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_2 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_2 <= _T_39; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_3 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_3 <= _T_41; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_4 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_4 <= _T_43; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_5 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_5 <= _T_45; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_6 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_6 <= _T_47; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_7 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_7 <= _T_49; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_8 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_8 <= _T_51; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_9 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_9 <= _T_53; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_10 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_10 <= _T_55; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_11 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_11 <= _T_57; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_12 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_12 <= _T_59; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_13 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_13 <= _T_61; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_14 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_14 <= _T_63; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_15 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_15 <= _T_65; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_16 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_16 <= _T_67; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_17 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_17 <= _T_69; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_18 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_18 <= _T_71; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_19 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_19 <= _T_73; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_20 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_20 <= _T_75; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_21 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_21 <= _T_77; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_22 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_22 <= _T_79; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_23 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_23 <= _T_81; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_24 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_24 <= _T_83; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_25 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_25 <= _T_85; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_26 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_26 <= _T_87; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_27 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_27 <= _T_89; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_28 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_28 <= _T_91; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_29 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_29 <= _T_93; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_30 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_30 <= _T_95; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 37:22]
      bits_31 <= 16'sh0; // @[VectorSerializer.scala 37:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      if (io_in_valid) begin // @[VectorSerializer.scala 55:23]
        bits_31 <= _T_97; // @[VectorSerializer.scala 56:12]
      end
    end
    if (reset) begin // @[VectorSerializer.scala 38:22]
      valid <= 1'h0; // @[VectorSerializer.scala 38:22]
    end else if (io_in_ready) begin // @[VectorSerializer.scala 54:21]
      valid <= io_in_valid;
    end
    if (reset) begin // @[Counter.scala 62:40]
      ctr <= 2'h0; // @[Counter.scala 62:40]
    end else if (_T) begin // @[Counter.scala 120:16]
      ctr <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bits_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  bits_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  bits_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  bits_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  bits_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  bits_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  bits_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  bits_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  bits_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  bits_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  bits_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  bits_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  bits_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  bits_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  bits_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  bits_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  bits_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  bits_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  bits_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  bits_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  bits_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  bits_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  bits_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  bits_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  bits_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  bits_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  bits_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  bits_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  bits_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  bits_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  bits_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  bits_31 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  ctr = _RAND_33[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DataCounter(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits,
  input          io_out_ready,
  output         io_out_valid,
  output [127:0] io_out_bits,
  output         io_len_ready,
  input          io_len_valid,
  input  [7:0]   io_len_bits
);
  wire  counter_clock; // @[Counter.scala 34:19]
  wire  counter_reset; // @[Counter.scala 34:19]
  wire  counter_io_value_ready; // @[Counter.scala 34:19]
  wire [7:0] counter_io_value_bits; // @[Counter.scala 34:19]
  wire  counter_io_resetValue; // @[Counter.scala 34:19]
  wire  _counter_io_resetValue_T = io_out_ready & io_out_valid; // @[Decoupled.scala 50:35]
  Counter_10 counter ( // @[Counter.scala 34:19]
    .clock(counter_clock),
    .reset(counter_reset),
    .io_value_ready(counter_io_value_ready),
    .io_value_bits(counter_io_value_bits),
    .io_resetValue(counter_io_resetValue)
  );
  assign io_in_ready = io_len_valid & io_out_ready; // @[DataCounter.scala 27:25]
  assign io_out_valid = io_in_valid & io_len_valid; // @[DataCounter.scala 26:28]
  assign io_out_bits = io_in_bits; // @[DataCounter.scala 25:15]
  assign io_len_ready = counter_io_value_bits == io_len_bits & (io_in_valid & io_out_ready); // @[DataCounter.scala 29:44 31:15 34:15]
  assign counter_clock = clock;
  assign counter_reset = reset;
  assign counter_io_value_ready = counter_io_value_bits == io_len_bits ? 1'h0 : _counter_io_resetValue_T; // @[DataCounter.scala 29:44 Counter.scala 36:22 DataCounter.scala 36:28]
  assign counter_io_resetValue = counter_io_value_bits == io_len_bits & _counter_io_resetValue_T; // @[DataCounter.scala 29:44 32:27 Counter.scala 35:21]
endmodule
module VectorDeserializer(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits,
  input          io_out_ready,
  output         io_out_valid,
  output [15:0]  io_out_bits_0,
  output [15:0]  io_out_bits_1,
  output [15:0]  io_out_bits_2,
  output [15:0]  io_out_bits_3,
  output [15:0]  io_out_bits_4,
  output [15:0]  io_out_bits_5,
  output [15:0]  io_out_bits_6,
  output [15:0]  io_out_bits_7,
  output [15:0]  io_out_bits_8,
  output [15:0]  io_out_bits_9,
  output [15:0]  io_out_bits_10,
  output [15:0]  io_out_bits_11,
  output [15:0]  io_out_bits_12,
  output [15:0]  io_out_bits_13,
  output [15:0]  io_out_bits_14,
  output [15:0]  io_out_bits_15,
  output [15:0]  io_out_bits_16,
  output [15:0]  io_out_bits_17,
  output [15:0]  io_out_bits_18,
  output [15:0]  io_out_bits_19,
  output [15:0]  io_out_bits_20,
  output [15:0]  io_out_bits_21,
  output [15:0]  io_out_bits_22,
  output [15:0]  io_out_bits_23,
  output [15:0]  io_out_bits_24,
  output [15:0]  io_out_bits_25,
  output [15:0]  io_out_bits_26,
  output [15:0]  io_out_bits_27,
  output [15:0]  io_out_bits_28,
  output [15:0]  io_out_bits_29,
  output [15:0]  io_out_bits_30,
  output [15:0]  io_out_bits_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] bits_0; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_1; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_2; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_3; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_4; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_5; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_6; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_7; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_8; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_9; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_10; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_11; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_12; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_13; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_14; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_15; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_16; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_17; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_18; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_19; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_20; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_21; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_22; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_23; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_24; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_25; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_26; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_27; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_28; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_29; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_30; // @[VectorDeserializer.scala 41:24]
  reg [15:0] bits_31; // @[VectorDeserializer.scala 41:24]
  reg  valid; // @[VectorDeserializer.scala 42:24]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
  reg [1:0] ctr; // @[Counter.scala 62:40]
  wire  wrap_wrap = ctr == 2'h3; // @[Counter.scala 74:24]
  wire [1:0] _wrap_value_T_1 = ctr + 2'h1; // @[Counter.scala 78:24]
  wire  wrap = _T & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire [5:0] _T_2 = ctr * 4'h8; // @[VectorDeserializer.scala 54:18]
  wire [6:0] _T_3 = {{1'd0}, _T_2}; // @[VectorDeserializer.scala 54:40]
  wire [15:0] _bits_T_65 = io_in_bits[15:0]; // @[VectorDeserializer.scala 37:57]
  wire [15:0] _GEN_2 = 5'h0 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_0); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_3 = 5'h1 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_1); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_4 = 5'h2 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_2); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_5 = 5'h3 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_3); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_6 = 5'h4 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_4); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_7 = 5'h5 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_5); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_8 = 5'h6 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_6); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_9 = 5'h7 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_7); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_10 = 5'h8 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_8); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_11 = 5'h9 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_9); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_12 = 5'ha == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_10); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_13 = 5'hb == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_11); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_14 = 5'hc == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_12); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_15 = 5'hd == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_13); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_16 = 5'he == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_14); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_17 = 5'hf == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_15); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_18 = 5'h10 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_16); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_19 = 5'h11 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_17); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_20 = 5'h12 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_18); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_21 = 5'h13 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_19); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_22 = 5'h14 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_20); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_23 = 5'h15 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_21); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_24 = 5'h16 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_22); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_25 = 5'h17 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_23); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_26 = 5'h18 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_24); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_27 = 5'h19 == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_25); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_28 = 5'h1a == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_26); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_29 = 5'h1b == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_27); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_30 = 5'h1c == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_28); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_31 = 5'h1d == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_29); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_32 = 5'h1e == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_30); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [15:0] _GEN_33 = 5'h1f == _T_3[4:0] ? $signed(_bits_T_65) : $signed(bits_31); // @[VectorDeserializer.scala 41:24 54:{47,47}]
  wire [5:0] _T_8 = _T_2 + 6'h1; // @[VectorDeserializer.scala 54:40]
  wire [15:0] _bits_T_67 = io_in_bits[31:16]; // @[VectorDeserializer.scala 37:57]
  wire [15:0] _GEN_34 = 5'h0 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_2); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_35 = 5'h1 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_3); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_36 = 5'h2 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_4); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_37 = 5'h3 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_5); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_38 = 5'h4 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_6); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_39 = 5'h5 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_7); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_40 = 5'h6 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_8); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_41 = 5'h7 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_9); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_42 = 5'h8 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_10); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_43 = 5'h9 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_11); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_44 = 5'ha == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_12); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_45 = 5'hb == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_13); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_46 = 5'hc == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_14); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_47 = 5'hd == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_15); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_48 = 5'he == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_16); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_49 = 5'hf == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_17); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_50 = 5'h10 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_18); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_51 = 5'h11 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_19); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_52 = 5'h12 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_20); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_53 = 5'h13 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_21); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_54 = 5'h14 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_22); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_55 = 5'h15 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_23); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_56 = 5'h16 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_24); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_57 = 5'h17 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_25); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_58 = 5'h18 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_26); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_59 = 5'h19 == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_27); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_60 = 5'h1a == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_28); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_61 = 5'h1b == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_29); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_62 = 5'h1c == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_30); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_63 = 5'h1d == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_31); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_64 = 5'h1e == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_32); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_65 = 5'h1f == _T_8[4:0] ? $signed(_bits_T_67) : $signed(_GEN_33); // @[VectorDeserializer.scala 54:{47,47}]
  wire [5:0] _T_12 = _T_2 + 6'h2; // @[VectorDeserializer.scala 54:40]
  wire [15:0] _bits_T_69 = io_in_bits[47:32]; // @[VectorDeserializer.scala 37:57]
  wire [15:0] _GEN_66 = 5'h0 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_34); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_67 = 5'h1 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_35); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_68 = 5'h2 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_36); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_69 = 5'h3 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_37); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_70 = 5'h4 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_38); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_71 = 5'h5 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_39); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_72 = 5'h6 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_40); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_73 = 5'h7 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_41); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_74 = 5'h8 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_42); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_75 = 5'h9 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_43); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_76 = 5'ha == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_44); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_77 = 5'hb == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_45); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_78 = 5'hc == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_46); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_79 = 5'hd == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_47); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_80 = 5'he == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_48); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_81 = 5'hf == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_49); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_82 = 5'h10 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_50); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_83 = 5'h11 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_51); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_84 = 5'h12 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_52); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_85 = 5'h13 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_53); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_86 = 5'h14 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_54); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_87 = 5'h15 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_55); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_88 = 5'h16 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_56); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_89 = 5'h17 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_57); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_90 = 5'h18 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_58); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_91 = 5'h19 == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_59); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_92 = 5'h1a == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_60); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_93 = 5'h1b == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_61); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_94 = 5'h1c == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_62); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_95 = 5'h1d == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_63); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_96 = 5'h1e == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_64); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_97 = 5'h1f == _T_12[4:0] ? $signed(_bits_T_69) : $signed(_GEN_65); // @[VectorDeserializer.scala 54:{47,47}]
  wire [5:0] _T_16 = _T_2 + 6'h3; // @[VectorDeserializer.scala 54:40]
  wire [15:0] _bits_T_71 = io_in_bits[63:48]; // @[VectorDeserializer.scala 37:57]
  wire [15:0] _GEN_98 = 5'h0 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_66); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_99 = 5'h1 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_67); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_100 = 5'h2 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_68); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_101 = 5'h3 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_69); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_102 = 5'h4 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_70); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_103 = 5'h5 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_71); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_104 = 5'h6 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_72); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_105 = 5'h7 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_73); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_106 = 5'h8 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_74); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_107 = 5'h9 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_75); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_108 = 5'ha == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_76); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_109 = 5'hb == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_77); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_110 = 5'hc == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_78); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_111 = 5'hd == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_79); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_112 = 5'he == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_80); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_113 = 5'hf == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_81); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_114 = 5'h10 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_82); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_115 = 5'h11 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_83); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_116 = 5'h12 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_84); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_117 = 5'h13 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_85); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_118 = 5'h14 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_86); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_119 = 5'h15 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_87); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_120 = 5'h16 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_88); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_121 = 5'h17 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_89); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_122 = 5'h18 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_90); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_123 = 5'h19 == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_91); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_124 = 5'h1a == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_92); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_125 = 5'h1b == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_93); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_126 = 5'h1c == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_94); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_127 = 5'h1d == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_95); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_128 = 5'h1e == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_96); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_129 = 5'h1f == _T_16[4:0] ? $signed(_bits_T_71) : $signed(_GEN_97); // @[VectorDeserializer.scala 54:{47,47}]
  wire [5:0] _T_20 = _T_2 + 6'h4; // @[VectorDeserializer.scala 54:40]
  wire [15:0] _bits_T_73 = io_in_bits[79:64]; // @[VectorDeserializer.scala 37:57]
  wire [15:0] _GEN_130 = 5'h0 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_98); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_131 = 5'h1 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_99); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_132 = 5'h2 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_100); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_133 = 5'h3 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_101); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_134 = 5'h4 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_102); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_135 = 5'h5 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_103); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_136 = 5'h6 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_104); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_137 = 5'h7 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_105); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_138 = 5'h8 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_106); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_139 = 5'h9 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_107); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_140 = 5'ha == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_108); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_141 = 5'hb == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_109); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_142 = 5'hc == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_110); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_143 = 5'hd == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_111); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_144 = 5'he == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_112); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_145 = 5'hf == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_113); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_146 = 5'h10 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_114); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_147 = 5'h11 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_115); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_148 = 5'h12 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_116); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_149 = 5'h13 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_117); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_150 = 5'h14 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_118); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_151 = 5'h15 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_119); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_152 = 5'h16 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_120); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_153 = 5'h17 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_121); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_154 = 5'h18 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_122); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_155 = 5'h19 == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_123); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_156 = 5'h1a == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_124); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_157 = 5'h1b == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_125); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_158 = 5'h1c == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_126); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_159 = 5'h1d == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_127); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_160 = 5'h1e == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_128); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_161 = 5'h1f == _T_20[4:0] ? $signed(_bits_T_73) : $signed(_GEN_129); // @[VectorDeserializer.scala 54:{47,47}]
  wire [5:0] _T_24 = _T_2 + 6'h5; // @[VectorDeserializer.scala 54:40]
  wire [15:0] _bits_T_75 = io_in_bits[95:80]; // @[VectorDeserializer.scala 37:57]
  wire [15:0] _GEN_162 = 5'h0 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_130); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_163 = 5'h1 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_131); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_164 = 5'h2 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_132); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_165 = 5'h3 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_133); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_166 = 5'h4 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_134); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_167 = 5'h5 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_135); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_168 = 5'h6 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_136); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_169 = 5'h7 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_137); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_170 = 5'h8 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_138); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_171 = 5'h9 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_139); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_172 = 5'ha == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_140); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_173 = 5'hb == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_141); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_174 = 5'hc == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_142); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_175 = 5'hd == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_143); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_176 = 5'he == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_144); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_177 = 5'hf == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_145); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_178 = 5'h10 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_146); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_179 = 5'h11 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_147); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_180 = 5'h12 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_148); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_181 = 5'h13 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_149); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_182 = 5'h14 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_150); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_183 = 5'h15 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_151); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_184 = 5'h16 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_152); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_185 = 5'h17 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_153); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_186 = 5'h18 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_154); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_187 = 5'h19 == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_155); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_188 = 5'h1a == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_156); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_189 = 5'h1b == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_157); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_190 = 5'h1c == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_158); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_191 = 5'h1d == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_159); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_192 = 5'h1e == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_160); // @[VectorDeserializer.scala 54:{47,47}]
  wire [15:0] _GEN_193 = 5'h1f == _T_24[4:0] ? $signed(_bits_T_75) : $signed(_GEN_161); // @[VectorDeserializer.scala 54:{47,47}]
  wire [5:0] _T_28 = _T_2 + 6'h6; // @[VectorDeserializer.scala 54:40]
  wire [15:0] _bits_T_77 = io_in_bits[111:96]; // @[VectorDeserializer.scala 37:57]
  wire [5:0] _T_32 = _T_2 + 6'h7; // @[VectorDeserializer.scala 54:40]
  wire [15:0] _bits_T_79 = io_in_bits[127:112]; // @[VectorDeserializer.scala 37:57]
  wire  _T_34 = io_out_ready & io_out_valid; // @[Decoupled.scala 50:35]
  assign io_in_ready = ~valid | io_out_ready; // @[VectorDeserializer.scala 50:27]
  assign io_out_valid = valid; // @[VectorDeserializer.scala 47:18]
  assign io_out_bits_0 = bits_0; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_1 = bits_1; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_2 = bits_2; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_3 = bits_3; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_4 = bits_4; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_5 = bits_5; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_6 = bits_6; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_7 = bits_7; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_8 = bits_8; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_9 = bits_9; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_10 = bits_10; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_11 = bits_11; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_12 = bits_12; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_13 = bits_13; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_14 = bits_14; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_15 = bits_15; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_16 = bits_16; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_17 = bits_17; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_18 = bits_18; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_19 = bits_19; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_20 = bits_20; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_21 = bits_21; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_22 = bits_22; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_23 = bits_23; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_24 = bits_24; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_25 = bits_25; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_26 = bits_26; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_27 = bits_27; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_28 = bits_28; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_29 = bits_29; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_30 = bits_30; // @[VectorDeserializer.scala 48:17]
  assign io_out_bits_31 = bits_31; // @[VectorDeserializer.scala 48:17]
  always @(posedge clock) begin
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_0 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h0 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_0 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h0 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_0 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_0 <= _GEN_162;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_1 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h1 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_1 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h1 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_1 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_1 <= _GEN_163;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_2 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h2 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_2 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h2 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_2 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_2 <= _GEN_164;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_3 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h3 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_3 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h3 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_3 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_3 <= _GEN_165;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_4 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h4 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_4 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h4 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_4 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_4 <= _GEN_166;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_5 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h5 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_5 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h5 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_5 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_5 <= _GEN_167;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_6 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h6 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_6 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h6 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_6 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_6 <= _GEN_168;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_7 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h7 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_7 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h7 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_7 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_7 <= _GEN_169;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_8 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h8 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_8 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h8 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_8 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_8 <= _GEN_170;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_9 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h9 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_9 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h9 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_9 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_9 <= _GEN_171;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_10 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'ha == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_10 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'ha == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_10 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_10 <= _GEN_172;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_11 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'hb == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_11 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'hb == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_11 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_11 <= _GEN_173;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_12 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'hc == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_12 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'hc == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_12 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_12 <= _GEN_174;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_13 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'hd == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_13 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'hd == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_13 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_13 <= _GEN_175;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_14 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'he == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_14 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'he == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_14 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_14 <= _GEN_176;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_15 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'hf == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_15 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'hf == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_15 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_15 <= _GEN_177;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_16 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h10 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_16 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h10 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_16 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_16 <= _GEN_178;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_17 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h11 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_17 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h11 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_17 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_17 <= _GEN_179;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_18 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h12 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_18 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h12 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_18 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_18 <= _GEN_180;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_19 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h13 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_19 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h13 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_19 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_19 <= _GEN_181;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_20 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h14 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_20 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h14 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_20 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_20 <= _GEN_182;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_21 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h15 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_21 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h15 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_21 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_21 <= _GEN_183;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_22 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h16 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_22 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h16 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_22 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_22 <= _GEN_184;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_23 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h17 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_23 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h17 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_23 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_23 <= _GEN_185;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_24 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h18 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_24 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h18 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_24 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_24 <= _GEN_186;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_25 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h19 == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_25 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h19 == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_25 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_25 <= _GEN_187;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_26 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h1a == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_26 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h1a == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_26 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_26 <= _GEN_188;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_27 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h1b == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_27 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h1b == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_27 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_27 <= _GEN_189;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_28 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h1c == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_28 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h1c == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_28 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_28 <= _GEN_190;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_29 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h1d == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_29 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h1d == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_29 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_29 <= _GEN_191;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_30 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h1e == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_30 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h1e == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_30 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_30 <= _GEN_192;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 41:24]
      bits_31 <= 16'sh0; // @[VectorDeserializer.scala 41:24]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      if (5'h1f == _T_32[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_31 <= _bits_T_79; // @[VectorDeserializer.scala 54:47]
      end else if (5'h1f == _T_28[4:0]) begin // @[VectorDeserializer.scala 54:47]
        bits_31 <= _bits_T_77; // @[VectorDeserializer.scala 54:47]
      end else begin
        bits_31 <= _GEN_193;
      end
    end
    if (reset) begin // @[VectorDeserializer.scala 42:24]
      valid <= 1'h0; // @[VectorDeserializer.scala 42:24]
    end else if (_T_34) begin // @[VectorDeserializer.scala 63:23]
      valid <= 1'h0; // @[VectorDeserializer.scala 64:13]
    end else if (_T) begin // @[VectorDeserializer.scala 52:22]
      valid <= wrap; // @[VectorDeserializer.scala 61:13]
    end
    if (reset) begin // @[Counter.scala 62:40]
      ctr <= 2'h0; // @[Counter.scala 62:40]
    end else if (_T) begin // @[Counter.scala 120:16]
      ctr <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bits_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  bits_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  bits_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  bits_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  bits_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  bits_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  bits_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  bits_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  bits_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  bits_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  bits_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  bits_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  bits_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  bits_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  bits_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  bits_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  bits_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  bits_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  bits_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  bits_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  bits_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  bits_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  bits_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  bits_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  bits_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  bits_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  bits_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  bits_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  bits_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  bits_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  bits_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  bits_31 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  ctr = _RAND_33[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Converter(
  input          clock,
  input          reset,
  output         io_mem_control_ready,
  input          io_mem_control_valid,
  input          io_mem_control_bits_write,
  input  [20:0]  io_mem_control_bits_address,
  input  [20:0]  io_mem_control_bits_size,
  input          io_mem_dataIn_ready,
  output         io_mem_dataIn_valid,
  output [15:0]  io_mem_dataIn_bits_0,
  output [15:0]  io_mem_dataIn_bits_1,
  output [15:0]  io_mem_dataIn_bits_2,
  output [15:0]  io_mem_dataIn_bits_3,
  output [15:0]  io_mem_dataIn_bits_4,
  output [15:0]  io_mem_dataIn_bits_5,
  output [15:0]  io_mem_dataIn_bits_6,
  output [15:0]  io_mem_dataIn_bits_7,
  output [15:0]  io_mem_dataIn_bits_8,
  output [15:0]  io_mem_dataIn_bits_9,
  output [15:0]  io_mem_dataIn_bits_10,
  output [15:0]  io_mem_dataIn_bits_11,
  output [15:0]  io_mem_dataIn_bits_12,
  output [15:0]  io_mem_dataIn_bits_13,
  output [15:0]  io_mem_dataIn_bits_14,
  output [15:0]  io_mem_dataIn_bits_15,
  output [15:0]  io_mem_dataIn_bits_16,
  output [15:0]  io_mem_dataIn_bits_17,
  output [15:0]  io_mem_dataIn_bits_18,
  output [15:0]  io_mem_dataIn_bits_19,
  output [15:0]  io_mem_dataIn_bits_20,
  output [15:0]  io_mem_dataIn_bits_21,
  output [15:0]  io_mem_dataIn_bits_22,
  output [15:0]  io_mem_dataIn_bits_23,
  output [15:0]  io_mem_dataIn_bits_24,
  output [15:0]  io_mem_dataIn_bits_25,
  output [15:0]  io_mem_dataIn_bits_26,
  output [15:0]  io_mem_dataIn_bits_27,
  output [15:0]  io_mem_dataIn_bits_28,
  output [15:0]  io_mem_dataIn_bits_29,
  output [15:0]  io_mem_dataIn_bits_30,
  output [15:0]  io_mem_dataIn_bits_31,
  output         io_mem_dataOut_ready,
  input          io_mem_dataOut_valid,
  input  [15:0]  io_mem_dataOut_bits_0,
  input  [15:0]  io_mem_dataOut_bits_1,
  input  [15:0]  io_mem_dataOut_bits_2,
  input  [15:0]  io_mem_dataOut_bits_3,
  input  [15:0]  io_mem_dataOut_bits_4,
  input  [15:0]  io_mem_dataOut_bits_5,
  input  [15:0]  io_mem_dataOut_bits_6,
  input  [15:0]  io_mem_dataOut_bits_7,
  input  [15:0]  io_mem_dataOut_bits_8,
  input  [15:0]  io_mem_dataOut_bits_9,
  input  [15:0]  io_mem_dataOut_bits_10,
  input  [15:0]  io_mem_dataOut_bits_11,
  input  [15:0]  io_mem_dataOut_bits_12,
  input  [15:0]  io_mem_dataOut_bits_13,
  input  [15:0]  io_mem_dataOut_bits_14,
  input  [15:0]  io_mem_dataOut_bits_15,
  input  [15:0]  io_mem_dataOut_bits_16,
  input  [15:0]  io_mem_dataOut_bits_17,
  input  [15:0]  io_mem_dataOut_bits_18,
  input  [15:0]  io_mem_dataOut_bits_19,
  input  [15:0]  io_mem_dataOut_bits_20,
  input  [15:0]  io_mem_dataOut_bits_21,
  input  [15:0]  io_mem_dataOut_bits_22,
  input  [15:0]  io_mem_dataOut_bits_23,
  input  [15:0]  io_mem_dataOut_bits_24,
  input  [15:0]  io_mem_dataOut_bits_25,
  input  [15:0]  io_mem_dataOut_bits_26,
  input  [15:0]  io_mem_dataOut_bits_27,
  input  [15:0]  io_mem_dataOut_bits_28,
  input  [15:0]  io_mem_dataOut_bits_29,
  input  [15:0]  io_mem_dataOut_bits_30,
  input  [15:0]  io_mem_dataOut_bits_31,
  input          io_axi_writeAddress_ready,
  output         io_axi_writeAddress_valid,
  output [31:0]  io_axi_writeAddress_bits_addr,
  output [7:0]   io_axi_writeAddress_bits_len,
  output [3:0]   io_axi_writeAddress_bits_cache,
  input          io_axi_writeData_ready,
  output         io_axi_writeData_valid,
  output [127:0] io_axi_writeData_bits_data,
  output         io_axi_writeResponse_ready,
  input          io_axi_writeResponse_valid,
  input          io_axi_readAddress_ready,
  output         io_axi_readAddress_valid,
  output [31:0]  io_axi_readAddress_bits_addr,
  output [7:0]   io_axi_readAddress_bits_len,
  output [3:0]   io_axi_readAddress_bits_cache,
  output         io_axi_readData_ready,
  input          io_axi_readData_valid,
  input  [127:0] io_axi_readData_bits_data,
  input          io_axi_readData_bits_last,
  input  [31:0]  io_addressOffset,
  input  [3:0]   io_cacheBehavior,
  input          io_timeout,
  input          io_tracepoint,
  input  [31:0]  io_programCounter
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  control_q_clock; // @[Converter.scala 65:25]
  wire  control_q_reset; // @[Converter.scala 65:25]
  wire  control_q_io_enq_ready; // @[Converter.scala 65:25]
  wire  control_q_io_enq_valid; // @[Converter.scala 65:25]
  wire  control_q_io_enq_bits_write; // @[Converter.scala 65:25]
  wire [20:0] control_q_io_enq_bits_address; // @[Converter.scala 65:25]
  wire [20:0] control_q_io_enq_bits_size; // @[Converter.scala 65:25]
  wire  control_q_io_deq_ready; // @[Converter.scala 65:25]
  wire  control_q_io_deq_valid; // @[Converter.scala 65:25]
  wire  control_q_io_deq_bits_write; // @[Converter.scala 65:25]
  wire [20:0] control_q_io_deq_bits_address; // @[Converter.scala 65:25]
  wire [20:0] control_q_io_deq_bits_size; // @[Converter.scala 65:25]
  wire  control_splitter_clock; // @[RequestSplitter.scala 69:26]
  wire  control_splitter_reset; // @[RequestSplitter.scala 69:26]
  wire  control_splitter_io_in_ready; // @[RequestSplitter.scala 69:26]
  wire  control_splitter_io_in_valid; // @[RequestSplitter.scala 69:26]
  wire  control_splitter_io_in_bits_write; // @[RequestSplitter.scala 69:26]
  wire [20:0] control_splitter_io_in_bits_address; // @[RequestSplitter.scala 69:26]
  wire [20:0] control_splitter_io_in_bits_size; // @[RequestSplitter.scala 69:26]
  wire  control_splitter_io_out_ready; // @[RequestSplitter.scala 69:26]
  wire  control_splitter_io_out_valid; // @[RequestSplitter.scala 69:26]
  wire  control_splitter_io_out_bits_write; // @[RequestSplitter.scala 69:26]
  wire [20:0] control_splitter_io_out_bits_address; // @[RequestSplitter.scala 69:26]
  wire [20:0] control_splitter_io_out_bits_size; // @[RequestSplitter.scala 69:26]
  wire  dataOut_clock; // @[Converter.scala 67:41]
  wire  dataOut_reset; // @[Converter.scala 67:41]
  wire  dataOut_io_enq_ready; // @[Converter.scala 67:41]
  wire  dataOut_io_enq_valid; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_0; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_1; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_2; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_3; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_4; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_5; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_6; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_7; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_8; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_9; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_10; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_11; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_12; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_13; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_14; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_15; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_16; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_17; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_18; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_19; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_20; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_21; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_22; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_23; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_24; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_25; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_26; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_27; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_28; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_29; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_30; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_enq_bits_31; // @[Converter.scala 67:41]
  wire  dataOut_io_deq_ready; // @[Converter.scala 67:41]
  wire  dataOut_io_deq_valid; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_0; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_1; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_2; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_3; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_4; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_5; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_6; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_7; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_8; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_9; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_10; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_11; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_12; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_13; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_14; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_15; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_16; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_17; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_18; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_19; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_20; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_21; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_22; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_23; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_24; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_25; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_26; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_27; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_28; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_29; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_30; // @[Converter.scala 67:41]
  wire [15:0] dataOut_io_deq_bits_31; // @[Converter.scala 67:41]
  wire  readData_clock; // @[Converter.scala 68:41]
  wire  readData_reset; // @[Converter.scala 68:41]
  wire  readData_io_enq_ready; // @[Converter.scala 68:41]
  wire  readData_io_enq_valid; // @[Converter.scala 68:41]
  wire [127:0] readData_io_enq_bits_data; // @[Converter.scala 68:41]
  wire  readData_io_enq_bits_last; // @[Converter.scala 68:41]
  wire  readData_io_deq_ready; // @[Converter.scala 68:41]
  wire  readData_io_deq_valid; // @[Converter.scala 68:41]
  wire [127:0] readData_io_deq_bits_data; // @[Converter.scala 68:41]
  wire  readData_io_deq_bits_last; // @[Converter.scala 68:41]
  wire  writeResponse_clock; // @[Converter.scala 69:41]
  wire  writeResponse_reset; // @[Converter.scala 69:41]
  wire  writeResponse_io_enq_ready; // @[Converter.scala 69:41]
  wire  writeResponse_io_enq_valid; // @[Converter.scala 69:41]
  wire  writeResponse_io_deq_ready; // @[Converter.scala 69:41]
  wire  writeResponse_io_deq_valid; // @[Converter.scala 69:41]
  wire  ser_clock; // @[Converter.scala 89:19]
  wire  ser_reset; // @[Converter.scala 89:19]
  wire  ser_io_in_ready; // @[Converter.scala 89:19]
  wire  ser_io_in_valid; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_0; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_1; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_2; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_3; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_4; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_5; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_6; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_7; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_8; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_9; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_10; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_11; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_12; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_13; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_14; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_15; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_16; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_17; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_18; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_19; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_20; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_21; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_22; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_23; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_24; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_25; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_26; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_27; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_28; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_29; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_30; // @[Converter.scala 89:19]
  wire [15:0] ser_io_in_bits_31; // @[Converter.scala 89:19]
  wire  ser_io_out_ready; // @[Converter.scala 89:19]
  wire  ser_io_out_valid; // @[Converter.scala 89:19]
  wire [127:0] ser_io_out_bits; // @[Converter.scala 89:19]
  wire  serCounter_clock; // @[Converter.scala 99:26]
  wire  serCounter_reset; // @[Converter.scala 99:26]
  wire  serCounter_io_in_ready; // @[Converter.scala 99:26]
  wire  serCounter_io_in_valid; // @[Converter.scala 99:26]
  wire [127:0] serCounter_io_in_bits; // @[Converter.scala 99:26]
  wire  serCounter_io_out_ready; // @[Converter.scala 99:26]
  wire  serCounter_io_out_valid; // @[Converter.scala 99:26]
  wire [127:0] serCounter_io_out_bits; // @[Converter.scala 99:26]
  wire  serCounter_io_len_ready; // @[Converter.scala 99:26]
  wire  serCounter_io_len_valid; // @[Converter.scala 99:26]
  wire [7:0] serCounter_io_len_bits; // @[Converter.scala 99:26]
  wire  des_clock; // @[Converter.scala 108:19]
  wire  des_reset; // @[Converter.scala 108:19]
  wire  des_io_in_ready; // @[Converter.scala 108:19]
  wire  des_io_in_valid; // @[Converter.scala 108:19]
  wire [127:0] des_io_in_bits; // @[Converter.scala 108:19]
  wire  des_io_out_ready; // @[Converter.scala 108:19]
  wire  des_io_out_valid; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_0; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_1; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_2; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_3; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_4; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_5; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_6; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_7; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_8; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_9; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_10; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_11; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_12; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_13; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_14; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_15; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_16; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_17; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_18; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_19; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_20; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_21; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_22; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_23; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_24; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_25; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_26; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_27; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_28; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_29; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_30; // @[Converter.scala 108:19]
  wire [15:0] des_io_out_bits_31; // @[Converter.scala 108:19]
  wire  writeEnqueue_clock; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueue_reset; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueue_io_in_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueue_io_in_valid; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueue_io_out_0_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueue_io_out_0_valid; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueue_io_out_1_ready; // @[MultiEnqueue.scala 182:43]
  wire  writeEnqueue_io_out_1_valid; // @[MultiEnqueue.scala 182:43]
  wire [27:0] address = control_splitter_io_out_bits_address * 7'h40; // @[Converter.scala 78:26]
  wire [20:0] _size_T_1 = control_splitter_io_out_bits_size + 21'h1; // @[Converter.scala 81:24]
  wire [23:0] _size_T_2 = _size_T_1 * 3'h4; // @[Converter.scala 81:31]
  wire [23:0] size = _size_T_2 - 24'h1; // @[Converter.scala 81:68]
  reg [7:0] writeResponseCount; // @[Converter.scala 123:35]
  reg [7:0] readResponseCount; // @[Converter.scala 124:35]
  wire  _canWrite_T_1 = writeResponseCount < 8'hff; // @[Converter.scala 126:56]
  wire  canWrite = readResponseCount == 8'h0 & writeResponseCount < 8'hff; // @[Converter.scala 126:33]
  wire  _canRead_T_1 = readResponseCount < 8'hff; // @[Converter.scala 128:56]
  wire  canRead = writeResponseCount == 8'h0 & readResponseCount < 8'hff; // @[Converter.scala 128:34]
  wire  writeRequested = io_axi_writeAddress_ready & io_axi_writeAddress_valid; // @[Converter.scala 129:50]
  wire  writeResponded = writeResponse_io_deq_ready & writeResponse_io_deq_valid; // @[Converter.scala 130:44]
  wire  readRequested = io_axi_readAddress_ready & io_axi_readAddress_valid; // @[Converter.scala 131:49]
  wire  readResponded = readData_io_deq_ready & readData_io_deq_valid & readData_io_deq_bits_last; // @[Converter.scala 132:57]
  wire [7:0] _writeResponseCount_T_1 = writeResponseCount + 8'h1; // @[Converter.scala 138:50]
  wire [7:0] _writeResponseCount_T_3 = writeResponseCount - 8'h1; // @[Converter.scala 143:48]
  wire [7:0] _readResponseCount_T_1 = readResponseCount + 8'h1; // @[Converter.scala 153:48]
  wire [7:0] _readResponseCount_T_3 = readResponseCount - 8'h1; // @[Converter.scala 158:46]
  wire [31:0] _GEN_15 = {{4'd0}, address}; // @[Converter.scala 168:15]
  Queue_36 control_q ( // @[Converter.scala 65:25]
    .clock(control_q_clock),
    .reset(control_q_reset),
    .io_enq_ready(control_q_io_enq_ready),
    .io_enq_valid(control_q_io_enq_valid),
    .io_enq_bits_write(control_q_io_enq_bits_write),
    .io_enq_bits_address(control_q_io_enq_bits_address),
    .io_enq_bits_size(control_q_io_enq_bits_size),
    .io_deq_ready(control_q_io_deq_ready),
    .io_deq_valid(control_q_io_deq_valid),
    .io_deq_bits_write(control_q_io_deq_bits_write),
    .io_deq_bits_address(control_q_io_deq_bits_address),
    .io_deq_bits_size(control_q_io_deq_bits_size)
  );
  RequestSplitter control_splitter ( // @[RequestSplitter.scala 69:26]
    .clock(control_splitter_clock),
    .reset(control_splitter_reset),
    .io_in_ready(control_splitter_io_in_ready),
    .io_in_valid(control_splitter_io_in_valid),
    .io_in_bits_write(control_splitter_io_in_bits_write),
    .io_in_bits_address(control_splitter_io_in_bits_address),
    .io_in_bits_size(control_splitter_io_in_bits_size),
    .io_out_ready(control_splitter_io_out_ready),
    .io_out_valid(control_splitter_io_out_valid),
    .io_out_bits_write(control_splitter_io_out_bits_write),
    .io_out_bits_address(control_splitter_io_out_bits_address),
    .io_out_bits_size(control_splitter_io_out_bits_size)
  );
  Queue_37 dataOut ( // @[Converter.scala 67:41]
    .clock(dataOut_clock),
    .reset(dataOut_reset),
    .io_enq_ready(dataOut_io_enq_ready),
    .io_enq_valid(dataOut_io_enq_valid),
    .io_enq_bits_0(dataOut_io_enq_bits_0),
    .io_enq_bits_1(dataOut_io_enq_bits_1),
    .io_enq_bits_2(dataOut_io_enq_bits_2),
    .io_enq_bits_3(dataOut_io_enq_bits_3),
    .io_enq_bits_4(dataOut_io_enq_bits_4),
    .io_enq_bits_5(dataOut_io_enq_bits_5),
    .io_enq_bits_6(dataOut_io_enq_bits_6),
    .io_enq_bits_7(dataOut_io_enq_bits_7),
    .io_enq_bits_8(dataOut_io_enq_bits_8),
    .io_enq_bits_9(dataOut_io_enq_bits_9),
    .io_enq_bits_10(dataOut_io_enq_bits_10),
    .io_enq_bits_11(dataOut_io_enq_bits_11),
    .io_enq_bits_12(dataOut_io_enq_bits_12),
    .io_enq_bits_13(dataOut_io_enq_bits_13),
    .io_enq_bits_14(dataOut_io_enq_bits_14),
    .io_enq_bits_15(dataOut_io_enq_bits_15),
    .io_enq_bits_16(dataOut_io_enq_bits_16),
    .io_enq_bits_17(dataOut_io_enq_bits_17),
    .io_enq_bits_18(dataOut_io_enq_bits_18),
    .io_enq_bits_19(dataOut_io_enq_bits_19),
    .io_enq_bits_20(dataOut_io_enq_bits_20),
    .io_enq_bits_21(dataOut_io_enq_bits_21),
    .io_enq_bits_22(dataOut_io_enq_bits_22),
    .io_enq_bits_23(dataOut_io_enq_bits_23),
    .io_enq_bits_24(dataOut_io_enq_bits_24),
    .io_enq_bits_25(dataOut_io_enq_bits_25),
    .io_enq_bits_26(dataOut_io_enq_bits_26),
    .io_enq_bits_27(dataOut_io_enq_bits_27),
    .io_enq_bits_28(dataOut_io_enq_bits_28),
    .io_enq_bits_29(dataOut_io_enq_bits_29),
    .io_enq_bits_30(dataOut_io_enq_bits_30),
    .io_enq_bits_31(dataOut_io_enq_bits_31),
    .io_deq_ready(dataOut_io_deq_ready),
    .io_deq_valid(dataOut_io_deq_valid),
    .io_deq_bits_0(dataOut_io_deq_bits_0),
    .io_deq_bits_1(dataOut_io_deq_bits_1),
    .io_deq_bits_2(dataOut_io_deq_bits_2),
    .io_deq_bits_3(dataOut_io_deq_bits_3),
    .io_deq_bits_4(dataOut_io_deq_bits_4),
    .io_deq_bits_5(dataOut_io_deq_bits_5),
    .io_deq_bits_6(dataOut_io_deq_bits_6),
    .io_deq_bits_7(dataOut_io_deq_bits_7),
    .io_deq_bits_8(dataOut_io_deq_bits_8),
    .io_deq_bits_9(dataOut_io_deq_bits_9),
    .io_deq_bits_10(dataOut_io_deq_bits_10),
    .io_deq_bits_11(dataOut_io_deq_bits_11),
    .io_deq_bits_12(dataOut_io_deq_bits_12),
    .io_deq_bits_13(dataOut_io_deq_bits_13),
    .io_deq_bits_14(dataOut_io_deq_bits_14),
    .io_deq_bits_15(dataOut_io_deq_bits_15),
    .io_deq_bits_16(dataOut_io_deq_bits_16),
    .io_deq_bits_17(dataOut_io_deq_bits_17),
    .io_deq_bits_18(dataOut_io_deq_bits_18),
    .io_deq_bits_19(dataOut_io_deq_bits_19),
    .io_deq_bits_20(dataOut_io_deq_bits_20),
    .io_deq_bits_21(dataOut_io_deq_bits_21),
    .io_deq_bits_22(dataOut_io_deq_bits_22),
    .io_deq_bits_23(dataOut_io_deq_bits_23),
    .io_deq_bits_24(dataOut_io_deq_bits_24),
    .io_deq_bits_25(dataOut_io_deq_bits_25),
    .io_deq_bits_26(dataOut_io_deq_bits_26),
    .io_deq_bits_27(dataOut_io_deq_bits_27),
    .io_deq_bits_28(dataOut_io_deq_bits_28),
    .io_deq_bits_29(dataOut_io_deq_bits_29),
    .io_deq_bits_30(dataOut_io_deq_bits_30),
    .io_deq_bits_31(dataOut_io_deq_bits_31)
  );
  Queue_38 readData ( // @[Converter.scala 68:41]
    .clock(readData_clock),
    .reset(readData_reset),
    .io_enq_ready(readData_io_enq_ready),
    .io_enq_valid(readData_io_enq_valid),
    .io_enq_bits_data(readData_io_enq_bits_data),
    .io_enq_bits_last(readData_io_enq_bits_last),
    .io_deq_ready(readData_io_deq_ready),
    .io_deq_valid(readData_io_deq_valid),
    .io_deq_bits_data(readData_io_deq_bits_data),
    .io_deq_bits_last(readData_io_deq_bits_last)
  );
  Queue_39 writeResponse ( // @[Converter.scala 69:41]
    .clock(writeResponse_clock),
    .reset(writeResponse_reset),
    .io_enq_ready(writeResponse_io_enq_ready),
    .io_enq_valid(writeResponse_io_enq_valid),
    .io_deq_ready(writeResponse_io_deq_ready),
    .io_deq_valid(writeResponse_io_deq_valid)
  );
  VectorSerializer ser ( // @[Converter.scala 89:19]
    .clock(ser_clock),
    .reset(ser_reset),
    .io_in_ready(ser_io_in_ready),
    .io_in_valid(ser_io_in_valid),
    .io_in_bits_0(ser_io_in_bits_0),
    .io_in_bits_1(ser_io_in_bits_1),
    .io_in_bits_2(ser_io_in_bits_2),
    .io_in_bits_3(ser_io_in_bits_3),
    .io_in_bits_4(ser_io_in_bits_4),
    .io_in_bits_5(ser_io_in_bits_5),
    .io_in_bits_6(ser_io_in_bits_6),
    .io_in_bits_7(ser_io_in_bits_7),
    .io_in_bits_8(ser_io_in_bits_8),
    .io_in_bits_9(ser_io_in_bits_9),
    .io_in_bits_10(ser_io_in_bits_10),
    .io_in_bits_11(ser_io_in_bits_11),
    .io_in_bits_12(ser_io_in_bits_12),
    .io_in_bits_13(ser_io_in_bits_13),
    .io_in_bits_14(ser_io_in_bits_14),
    .io_in_bits_15(ser_io_in_bits_15),
    .io_in_bits_16(ser_io_in_bits_16),
    .io_in_bits_17(ser_io_in_bits_17),
    .io_in_bits_18(ser_io_in_bits_18),
    .io_in_bits_19(ser_io_in_bits_19),
    .io_in_bits_20(ser_io_in_bits_20),
    .io_in_bits_21(ser_io_in_bits_21),
    .io_in_bits_22(ser_io_in_bits_22),
    .io_in_bits_23(ser_io_in_bits_23),
    .io_in_bits_24(ser_io_in_bits_24),
    .io_in_bits_25(ser_io_in_bits_25),
    .io_in_bits_26(ser_io_in_bits_26),
    .io_in_bits_27(ser_io_in_bits_27),
    .io_in_bits_28(ser_io_in_bits_28),
    .io_in_bits_29(ser_io_in_bits_29),
    .io_in_bits_30(ser_io_in_bits_30),
    .io_in_bits_31(ser_io_in_bits_31),
    .io_out_ready(ser_io_out_ready),
    .io_out_valid(ser_io_out_valid),
    .io_out_bits(ser_io_out_bits)
  );
  DataCounter serCounter ( // @[Converter.scala 99:26]
    .clock(serCounter_clock),
    .reset(serCounter_reset),
    .io_in_ready(serCounter_io_in_ready),
    .io_in_valid(serCounter_io_in_valid),
    .io_in_bits(serCounter_io_in_bits),
    .io_out_ready(serCounter_io_out_ready),
    .io_out_valid(serCounter_io_out_valid),
    .io_out_bits(serCounter_io_out_bits),
    .io_len_ready(serCounter_io_len_ready),
    .io_len_valid(serCounter_io_len_valid),
    .io_len_bits(serCounter_io_len_bits)
  );
  VectorDeserializer des ( // @[Converter.scala 108:19]
    .clock(des_clock),
    .reset(des_reset),
    .io_in_ready(des_io_in_ready),
    .io_in_valid(des_io_in_valid),
    .io_in_bits(des_io_in_bits),
    .io_out_ready(des_io_out_ready),
    .io_out_valid(des_io_out_valid),
    .io_out_bits_0(des_io_out_bits_0),
    .io_out_bits_1(des_io_out_bits_1),
    .io_out_bits_2(des_io_out_bits_2),
    .io_out_bits_3(des_io_out_bits_3),
    .io_out_bits_4(des_io_out_bits_4),
    .io_out_bits_5(des_io_out_bits_5),
    .io_out_bits_6(des_io_out_bits_6),
    .io_out_bits_7(des_io_out_bits_7),
    .io_out_bits_8(des_io_out_bits_8),
    .io_out_bits_9(des_io_out_bits_9),
    .io_out_bits_10(des_io_out_bits_10),
    .io_out_bits_11(des_io_out_bits_11),
    .io_out_bits_12(des_io_out_bits_12),
    .io_out_bits_13(des_io_out_bits_13),
    .io_out_bits_14(des_io_out_bits_14),
    .io_out_bits_15(des_io_out_bits_15),
    .io_out_bits_16(des_io_out_bits_16),
    .io_out_bits_17(des_io_out_bits_17),
    .io_out_bits_18(des_io_out_bits_18),
    .io_out_bits_19(des_io_out_bits_19),
    .io_out_bits_20(des_io_out_bits_20),
    .io_out_bits_21(des_io_out_bits_21),
    .io_out_bits_22(des_io_out_bits_22),
    .io_out_bits_23(des_io_out_bits_23),
    .io_out_bits_24(des_io_out_bits_24),
    .io_out_bits_25(des_io_out_bits_25),
    .io_out_bits_26(des_io_out_bits_26),
    .io_out_bits_27(des_io_out_bits_27),
    .io_out_bits_28(des_io_out_bits_28),
    .io_out_bits_29(des_io_out_bits_29),
    .io_out_bits_30(des_io_out_bits_30),
    .io_out_bits_31(des_io_out_bits_31)
  );
  MultiEnqueue_1 writeEnqueue ( // @[MultiEnqueue.scala 182:43]
    .clock(writeEnqueue_clock),
    .reset(writeEnqueue_reset),
    .io_in_ready(writeEnqueue_io_in_ready),
    .io_in_valid(writeEnqueue_io_in_valid),
    .io_out_0_ready(writeEnqueue_io_out_0_ready),
    .io_out_0_valid(writeEnqueue_io_out_0_valid),
    .io_out_1_ready(writeEnqueue_io_out_1_ready),
    .io_out_1_valid(writeEnqueue_io_out_1_valid)
  );
  assign io_mem_control_ready = control_q_io_enq_ready; // @[Converter.scala 65:25]
  assign io_mem_dataIn_valid = des_io_out_valid; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_0 = des_io_out_bits_0; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_1 = des_io_out_bits_1; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_2 = des_io_out_bits_2; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_3 = des_io_out_bits_3; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_4 = des_io_out_bits_4; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_5 = des_io_out_bits_5; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_6 = des_io_out_bits_6; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_7 = des_io_out_bits_7; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_8 = des_io_out_bits_8; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_9 = des_io_out_bits_9; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_10 = des_io_out_bits_10; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_11 = des_io_out_bits_11; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_12 = des_io_out_bits_12; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_13 = des_io_out_bits_13; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_14 = des_io_out_bits_14; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_15 = des_io_out_bits_15; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_16 = des_io_out_bits_16; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_17 = des_io_out_bits_17; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_18 = des_io_out_bits_18; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_19 = des_io_out_bits_19; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_20 = des_io_out_bits_20; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_21 = des_io_out_bits_21; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_22 = des_io_out_bits_22; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_23 = des_io_out_bits_23; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_24 = des_io_out_bits_24; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_25 = des_io_out_bits_25; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_26 = des_io_out_bits_26; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_27 = des_io_out_bits_27; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_28 = des_io_out_bits_28; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_29 = des_io_out_bits_29; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_30 = des_io_out_bits_30; // @[Converter.scala 116:17]
  assign io_mem_dataIn_bits_31 = des_io_out_bits_31; // @[Converter.scala 116:17]
  assign io_mem_dataOut_ready = dataOut_io_enq_ready; // @[Converter.scala 67:41]
  assign io_axi_writeAddress_valid = control_splitter_io_out_bits_write & writeEnqueue_io_out_0_valid; // @[Converter.scala 207:28 172:29 212:31]
  assign io_axi_writeAddress_bits_addr = _GEN_15 + io_addressOffset; // @[Converter.scala 168:15]
  assign io_axi_writeAddress_bits_len = size[7:0]; // @[Address.scala 28:9]
  assign io_axi_writeAddress_bits_cache = io_cacheBehavior; // @[Address.scala 30:34]
  assign io_axi_writeData_valid = serCounter_io_out_valid; // @[Converter.scala 179:26]
  assign io_axi_writeData_bits_data = serCounter_io_out_bits; // @[WriteData.scala 20:15]
  assign io_axi_writeResponse_ready = writeResponse_io_enq_ready; // @[Converter.scala 69:41]
  assign io_axi_readAddress_valid = control_splitter_io_out_bits_write ? 1'h0 : control_splitter_io_out_valid & canRead; // @[Converter.scala 194:28 207:28 216:30]
  assign io_axi_readAddress_bits_addr = _GEN_15 + io_addressOffset; // @[Converter.scala 190:15]
  assign io_axi_readAddress_bits_len = size[7:0]; // @[Address.scala 28:9]
  assign io_axi_readAddress_bits_cache = io_cacheBehavior; // @[Address.scala 30:34]
  assign io_axi_readData_ready = readData_io_enq_ready; // @[Converter.scala 68:41]
  assign control_q_clock = clock;
  assign control_q_reset = reset;
  assign control_q_io_enq_valid = io_mem_control_valid; // @[Converter.scala 65:25]
  assign control_q_io_enq_bits_write = io_mem_control_bits_write; // @[Converter.scala 65:25]
  assign control_q_io_enq_bits_address = io_mem_control_bits_address; // @[Converter.scala 65:25]
  assign control_q_io_enq_bits_size = io_mem_control_bits_size; // @[Converter.scala 65:25]
  assign control_q_io_deq_ready = control_splitter_io_in_ready; // @[RequestSplitter.scala 70:20]
  assign control_splitter_clock = clock;
  assign control_splitter_reset = reset;
  assign control_splitter_io_in_valid = control_q_io_deq_valid; // @[RequestSplitter.scala 70:20]
  assign control_splitter_io_in_bits_write = control_q_io_deq_bits_write; // @[RequestSplitter.scala 70:20]
  assign control_splitter_io_in_bits_address = control_q_io_deq_bits_address; // @[RequestSplitter.scala 70:20]
  assign control_splitter_io_in_bits_size = control_q_io_deq_bits_size; // @[RequestSplitter.scala 70:20]
  assign control_splitter_io_out_ready = control_splitter_io_out_bits_write ? writeEnqueue_io_in_ready :
    io_axi_readAddress_ready & canRead; // @[Converter.scala 207:28 209:19 217:19]
  assign dataOut_clock = clock;
  assign dataOut_reset = reset;
  assign dataOut_io_enq_valid = io_mem_dataOut_valid; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_0 = io_mem_dataOut_bits_0; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_1 = io_mem_dataOut_bits_1; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_2 = io_mem_dataOut_bits_2; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_3 = io_mem_dataOut_bits_3; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_4 = io_mem_dataOut_bits_4; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_5 = io_mem_dataOut_bits_5; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_6 = io_mem_dataOut_bits_6; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_7 = io_mem_dataOut_bits_7; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_8 = io_mem_dataOut_bits_8; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_9 = io_mem_dataOut_bits_9; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_10 = io_mem_dataOut_bits_10; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_11 = io_mem_dataOut_bits_11; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_12 = io_mem_dataOut_bits_12; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_13 = io_mem_dataOut_bits_13; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_14 = io_mem_dataOut_bits_14; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_15 = io_mem_dataOut_bits_15; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_16 = io_mem_dataOut_bits_16; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_17 = io_mem_dataOut_bits_17; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_18 = io_mem_dataOut_bits_18; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_19 = io_mem_dataOut_bits_19; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_20 = io_mem_dataOut_bits_20; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_21 = io_mem_dataOut_bits_21; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_22 = io_mem_dataOut_bits_22; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_23 = io_mem_dataOut_bits_23; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_24 = io_mem_dataOut_bits_24; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_25 = io_mem_dataOut_bits_25; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_26 = io_mem_dataOut_bits_26; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_27 = io_mem_dataOut_bits_27; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_28 = io_mem_dataOut_bits_28; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_29 = io_mem_dataOut_bits_29; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_30 = io_mem_dataOut_bits_30; // @[Converter.scala 67:41]
  assign dataOut_io_enq_bits_31 = io_mem_dataOut_bits_31; // @[Converter.scala 67:41]
  assign dataOut_io_deq_ready = ser_io_in_ready; // @[Converter.scala 97:13]
  assign readData_clock = clock;
  assign readData_reset = reset;
  assign readData_io_enq_valid = io_axi_readData_valid; // @[Converter.scala 68:41]
  assign readData_io_enq_bits_data = io_axi_readData_bits_data; // @[Converter.scala 68:41]
  assign readData_io_enq_bits_last = io_axi_readData_bits_last; // @[Converter.scala 68:41]
  assign readData_io_deq_ready = des_io_in_ready; // @[Converter.scala 201:18]
  assign writeResponse_clock = clock;
  assign writeResponse_reset = reset;
  assign writeResponse_io_enq_valid = io_axi_writeResponse_valid; // @[Converter.scala 69:41]
  assign writeResponse_io_deq_ready = 1'h1; // @[Converter.scala 184:23]
  assign ser_clock = clock;
  assign ser_reset = reset;
  assign ser_io_in_valid = dataOut_io_deq_valid; // @[Converter.scala 97:13]
  assign ser_io_in_bits_0 = dataOut_io_deq_bits_0; // @[Converter.scala 97:13]
  assign ser_io_in_bits_1 = dataOut_io_deq_bits_1; // @[Converter.scala 97:13]
  assign ser_io_in_bits_2 = dataOut_io_deq_bits_2; // @[Converter.scala 97:13]
  assign ser_io_in_bits_3 = dataOut_io_deq_bits_3; // @[Converter.scala 97:13]
  assign ser_io_in_bits_4 = dataOut_io_deq_bits_4; // @[Converter.scala 97:13]
  assign ser_io_in_bits_5 = dataOut_io_deq_bits_5; // @[Converter.scala 97:13]
  assign ser_io_in_bits_6 = dataOut_io_deq_bits_6; // @[Converter.scala 97:13]
  assign ser_io_in_bits_7 = dataOut_io_deq_bits_7; // @[Converter.scala 97:13]
  assign ser_io_in_bits_8 = dataOut_io_deq_bits_8; // @[Converter.scala 97:13]
  assign ser_io_in_bits_9 = dataOut_io_deq_bits_9; // @[Converter.scala 97:13]
  assign ser_io_in_bits_10 = dataOut_io_deq_bits_10; // @[Converter.scala 97:13]
  assign ser_io_in_bits_11 = dataOut_io_deq_bits_11; // @[Converter.scala 97:13]
  assign ser_io_in_bits_12 = dataOut_io_deq_bits_12; // @[Converter.scala 97:13]
  assign ser_io_in_bits_13 = dataOut_io_deq_bits_13; // @[Converter.scala 97:13]
  assign ser_io_in_bits_14 = dataOut_io_deq_bits_14; // @[Converter.scala 97:13]
  assign ser_io_in_bits_15 = dataOut_io_deq_bits_15; // @[Converter.scala 97:13]
  assign ser_io_in_bits_16 = dataOut_io_deq_bits_16; // @[Converter.scala 97:13]
  assign ser_io_in_bits_17 = dataOut_io_deq_bits_17; // @[Converter.scala 97:13]
  assign ser_io_in_bits_18 = dataOut_io_deq_bits_18; // @[Converter.scala 97:13]
  assign ser_io_in_bits_19 = dataOut_io_deq_bits_19; // @[Converter.scala 97:13]
  assign ser_io_in_bits_20 = dataOut_io_deq_bits_20; // @[Converter.scala 97:13]
  assign ser_io_in_bits_21 = dataOut_io_deq_bits_21; // @[Converter.scala 97:13]
  assign ser_io_in_bits_22 = dataOut_io_deq_bits_22; // @[Converter.scala 97:13]
  assign ser_io_in_bits_23 = dataOut_io_deq_bits_23; // @[Converter.scala 97:13]
  assign ser_io_in_bits_24 = dataOut_io_deq_bits_24; // @[Converter.scala 97:13]
  assign ser_io_in_bits_25 = dataOut_io_deq_bits_25; // @[Converter.scala 97:13]
  assign ser_io_in_bits_26 = dataOut_io_deq_bits_26; // @[Converter.scala 97:13]
  assign ser_io_in_bits_27 = dataOut_io_deq_bits_27; // @[Converter.scala 97:13]
  assign ser_io_in_bits_28 = dataOut_io_deq_bits_28; // @[Converter.scala 97:13]
  assign ser_io_in_bits_29 = dataOut_io_deq_bits_29; // @[Converter.scala 97:13]
  assign ser_io_in_bits_30 = dataOut_io_deq_bits_30; // @[Converter.scala 97:13]
  assign ser_io_in_bits_31 = dataOut_io_deq_bits_31; // @[Converter.scala 97:13]
  assign ser_io_out_ready = serCounter_io_in_ready; // @[Converter.scala 102:20]
  assign serCounter_clock = clock;
  assign serCounter_reset = reset;
  assign serCounter_io_in_valid = ser_io_out_valid; // @[Converter.scala 102:20]
  assign serCounter_io_in_bits = ser_io_out_bits; // @[Converter.scala 102:20]
  assign serCounter_io_out_ready = io_axi_writeData_ready; // @[Converter.scala 180:16]
  assign serCounter_io_len_valid = control_splitter_io_out_bits_write & writeEnqueue_io_out_1_valid; // @[Converter.scala 104:27 207:28 214:29]
  assign serCounter_io_len_bits = size[7:0]; // @[Converter.scala 103:26]
  assign des_clock = clock;
  assign des_reset = reset;
  assign des_io_in_valid = readData_io_deq_valid; // @[Converter.scala 200:19]
  assign des_io_in_bits = readData_io_deq_bits_data; // @[Converter.scala 199:18]
  assign des_io_out_ready = io_mem_dataIn_ready; // @[Converter.scala 116:17]
  assign writeEnqueue_clock = clock;
  assign writeEnqueue_reset = reset;
  assign writeEnqueue_io_in_valid = control_splitter_io_out_bits_write & (control_splitter_io_out_valid & canWrite); // @[Converter.scala 207:28 208:30 MultiEnqueue.scala 40:17]
  assign writeEnqueue_io_out_0_ready = control_splitter_io_out_bits_write & io_axi_writeAddress_ready; // @[Converter.scala 207:28 211:34 MultiEnqueue.scala 42:18]
  assign writeEnqueue_io_out_1_ready = control_splitter_io_out_bits_write & serCounter_io_len_ready; // @[Converter.scala 207:28 213:34 MultiEnqueue.scala 42:18]
  always @(posedge clock) begin
    if (reset) begin // @[Converter.scala 123:35]
      writeResponseCount <= 8'h0; // @[Converter.scala 123:35]
    end else if (writeRequested) begin // @[Converter.scala 133:24]
      if (!(writeResponded)) begin // @[Converter.scala 134:26]
        if (_canWrite_T_1) begin // @[Converter.scala 137:62]
          writeResponseCount <= _writeResponseCount_T_1; // @[Converter.scala 138:28]
        end
      end
    end else if (writeResponded & writeResponseCount > 8'h0) begin // @[Converter.scala 142:54]
      writeResponseCount <= _writeResponseCount_T_3; // @[Converter.scala 143:26]
    end
    if (reset) begin // @[Converter.scala 124:35]
      readResponseCount <= 8'h0; // @[Converter.scala 124:35]
    end else if (readRequested) begin // @[Converter.scala 148:23]
      if (!(readResponded)) begin // @[Converter.scala 149:25]
        if (_canRead_T_1) begin // @[Converter.scala 152:61]
          readResponseCount <= _readResponseCount_T_1; // @[Converter.scala 153:27]
        end
      end
    end else if (readResponded & readResponseCount > 8'h0) begin // @[Converter.scala 157:52]
      readResponseCount <= _readResponseCount_T_3; // @[Converter.scala 158:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeResponseCount = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  readResponseCount = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_40(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [3:0]  io_enq_bits_cache,
  input         io_deq_ready,
  output        io_deq_valid,
  output [5:0]  io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output [1:0]  io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] ram_id [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [5:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_addr [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_addr_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_len [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_burst [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_lock [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_lock_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_lock_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_lock_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_lock_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_lock_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_lock_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_cache [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_cache_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_cache_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_cache_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_prot [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_prot_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_prot_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_prot_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_qos [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_qos_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_qos_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_qos_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_qos_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_qos_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_qos_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = value_1;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_id_MPORT_data = 6'h0;
  assign ram_id_MPORT_addr = value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = value_1;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = value_1;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = 3'h4;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = value_1;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_burst_MPORT_data = 2'h1;
  assign ram_burst_MPORT_addr = value;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_lock_io_deq_bits_MPORT_en = 1'h1;
  assign ram_lock_io_deq_bits_MPORT_addr = value_1;
  assign ram_lock_io_deq_bits_MPORT_data = ram_lock[ram_lock_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_lock_MPORT_data = 2'h0;
  assign ram_lock_MPORT_addr = value;
  assign ram_lock_MPORT_mask = 1'h1;
  assign ram_lock_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_cache_io_deq_bits_MPORT_en = 1'h1;
  assign ram_cache_io_deq_bits_MPORT_addr = value_1;
  assign ram_cache_io_deq_bits_MPORT_data = ram_cache[ram_cache_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_cache_MPORT_data = io_enq_bits_cache;
  assign ram_cache_MPORT_addr = value;
  assign ram_cache_MPORT_mask = 1'h1;
  assign ram_cache_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_prot_io_deq_bits_MPORT_en = 1'h1;
  assign ram_prot_io_deq_bits_MPORT_addr = value_1;
  assign ram_prot_io_deq_bits_MPORT_data = ram_prot[ram_prot_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_prot_MPORT_data = 3'h0;
  assign ram_prot_MPORT_addr = value;
  assign ram_prot_MPORT_mask = 1'h1;
  assign ram_prot_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qos_io_deq_bits_MPORT_en = 1'h1;
  assign ram_qos_io_deq_bits_MPORT_addr = value_1;
  assign ram_qos_io_deq_bits_MPORT_data = ram_qos[ram_qos_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_qos_MPORT_data = 4'h0;
  assign ram_qos_MPORT_addr = value;
  assign ram_qos_MPORT_mask = 1'h1;
  assign ram_qos_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_burst = ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_lock = ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_cache = ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_prot = ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_qos = ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_lock_MPORT_en & ram_lock_MPORT_mask) begin
      ram_lock[ram_lock_MPORT_addr] <= ram_lock_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_cache_MPORT_en & ram_cache_MPORT_mask) begin
      ram_cache[ram_cache_MPORT_addr] <= ram_cache_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_prot_MPORT_en & ram_prot_MPORT_mask) begin
      ram_prot[ram_prot_MPORT_addr] <= ram_prot_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_qos_MPORT_en & ram_qos_MPORT_mask) begin
      ram_qos[ram_qos_MPORT_addr] <= ram_qos_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      value <= value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      value_1 <= value_1 + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_lock[initvar] = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_cache[initvar] = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_prot[initvar] = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_qos[initvar] = _RAND_8[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  value = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  value_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  maybe_full = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_42(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits_data,
  input          io_deq_ready,
  output         io_deq_valid,
  output [5:0]   io_deq_bits_id,
  output [127:0] io_deq_bits_data,
  output [15:0]  io_deq_bits_strb
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] ram_id [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [5:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg [127:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [127:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [127:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg [15:0] ram_strb [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_strb_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [15:0] ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [15:0] ram_strb_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_strb_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_strb_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_strb_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = value_1;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_id_MPORT_data = 6'h0;
  assign ram_id_MPORT_addr = value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_strb_io_deq_bits_MPORT_en = 1'h1;
  assign ram_strb_io_deq_bits_MPORT_addr = value_1;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_strb_MPORT_data = 16'hffff;
  assign ram_strb_MPORT_addr = value;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_strb = ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      value <= value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      value_1 <= value_1 + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[5:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[127:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_strb[initvar] = _RAND_2[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_45(
  input          clock,
  input          reset,
  output         io_in_writeAddress_ready,
  input          io_in_writeAddress_valid,
  input  [31:0]  io_in_writeAddress_bits_addr,
  input  [7:0]   io_in_writeAddress_bits_len,
  input  [3:0]   io_in_writeAddress_bits_cache,
  output         io_in_writeData_ready,
  input          io_in_writeData_valid,
  input  [127:0] io_in_writeData_bits_data,
  input          io_in_writeResponse_ready,
  output         io_in_writeResponse_valid,
  output         io_in_readAddress_ready,
  input          io_in_readAddress_valid,
  input  [31:0]  io_in_readAddress_bits_addr,
  input  [7:0]   io_in_readAddress_bits_len,
  input  [3:0]   io_in_readAddress_bits_cache,
  input          io_in_readData_ready,
  output         io_in_readData_valid,
  output [127:0] io_in_readData_bits_data,
  output         io_in_readData_bits_last,
  input          io_out_writeAddress_ready,
  output         io_out_writeAddress_valid,
  output [5:0]   io_out_writeAddress_bits_id,
  output [31:0]  io_out_writeAddress_bits_addr,
  output [7:0]   io_out_writeAddress_bits_len,
  output [2:0]   io_out_writeAddress_bits_size,
  output [1:0]   io_out_writeAddress_bits_burst,
  output [1:0]   io_out_writeAddress_bits_lock,
  output [3:0]   io_out_writeAddress_bits_cache,
  output [2:0]   io_out_writeAddress_bits_prot,
  output [3:0]   io_out_writeAddress_bits_qos,
  input          io_out_writeData_ready,
  output         io_out_writeData_valid,
  output [5:0]   io_out_writeData_bits_id,
  output [127:0] io_out_writeData_bits_data,
  output [15:0]  io_out_writeData_bits_strb,
  output         io_out_writeResponse_ready,
  input          io_out_writeResponse_valid,
  input          io_out_readAddress_ready,
  output         io_out_readAddress_valid,
  output [5:0]   io_out_readAddress_bits_id,
  output [31:0]  io_out_readAddress_bits_addr,
  output [7:0]   io_out_readAddress_bits_len,
  output [2:0]   io_out_readAddress_bits_size,
  output [1:0]   io_out_readAddress_bits_burst,
  output [1:0]   io_out_readAddress_bits_lock,
  output [3:0]   io_out_readAddress_bits_cache,
  output [2:0]   io_out_readAddress_bits_prot,
  output [3:0]   io_out_readAddress_bits_qos,
  output         io_out_readData_ready,
  input          io_out_readData_valid,
  input  [127:0] io_out_readData_bits_data,
  input          io_out_readData_bits_last
);
  wire  io_out_readAddress_q_clock; // @[Decoupled.scala 361:21]
  wire  io_out_readAddress_q_reset; // @[Decoupled.scala 361:21]
  wire  io_out_readAddress_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_readAddress_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] io_out_readAddress_q_io_enq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] io_out_readAddress_q_io_enq_bits_len; // @[Decoupled.scala 361:21]
  wire [3:0] io_out_readAddress_q_io_enq_bits_cache; // @[Decoupled.scala 361:21]
  wire  io_out_readAddress_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_readAddress_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [5:0] io_out_readAddress_q_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] io_out_readAddress_q_io_deq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] io_out_readAddress_q_io_deq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_readAddress_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] io_out_readAddress_q_io_deq_bits_burst; // @[Decoupled.scala 361:21]
  wire [1:0] io_out_readAddress_q_io_deq_bits_lock; // @[Decoupled.scala 361:21]
  wire [3:0] io_out_readAddress_q_io_deq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_readAddress_q_io_deq_bits_prot; // @[Decoupled.scala 361:21]
  wire [3:0] io_out_readAddress_q_io_deq_bits_qos; // @[Decoupled.scala 361:21]
  wire  io_out_writeAddress_q_clock; // @[Decoupled.scala 361:21]
  wire  io_out_writeAddress_q_reset; // @[Decoupled.scala 361:21]
  wire  io_out_writeAddress_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_writeAddress_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] io_out_writeAddress_q_io_enq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] io_out_writeAddress_q_io_enq_bits_len; // @[Decoupled.scala 361:21]
  wire [3:0] io_out_writeAddress_q_io_enq_bits_cache; // @[Decoupled.scala 361:21]
  wire  io_out_writeAddress_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_writeAddress_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [5:0] io_out_writeAddress_q_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] io_out_writeAddress_q_io_deq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] io_out_writeAddress_q_io_deq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_writeAddress_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] io_out_writeAddress_q_io_deq_bits_burst; // @[Decoupled.scala 361:21]
  wire [1:0] io_out_writeAddress_q_io_deq_bits_lock; // @[Decoupled.scala 361:21]
  wire [3:0] io_out_writeAddress_q_io_deq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_writeAddress_q_io_deq_bits_prot; // @[Decoupled.scala 361:21]
  wire [3:0] io_out_writeAddress_q_io_deq_bits_qos; // @[Decoupled.scala 361:21]
  wire  io_out_writeData_q_clock; // @[Decoupled.scala 361:21]
  wire  io_out_writeData_q_reset; // @[Decoupled.scala 361:21]
  wire  io_out_writeData_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_writeData_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [127:0] io_out_writeData_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  io_out_writeData_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_writeData_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [5:0] io_out_writeData_q_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [127:0] io_out_writeData_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [15:0] io_out_writeData_q_io_deq_bits_strb; // @[Decoupled.scala 361:21]
  wire  io_in_readData_q_clock; // @[Decoupled.scala 361:21]
  wire  io_in_readData_q_reset; // @[Decoupled.scala 361:21]
  wire  io_in_readData_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  io_in_readData_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [127:0] io_in_readData_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  io_in_readData_q_io_enq_bits_last; // @[Decoupled.scala 361:21]
  wire  io_in_readData_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  io_in_readData_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [127:0] io_in_readData_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire  io_in_readData_q_io_deq_bits_last; // @[Decoupled.scala 361:21]
  wire  io_in_writeResponse_q_clock; // @[Decoupled.scala 361:21]
  wire  io_in_writeResponse_q_reset; // @[Decoupled.scala 361:21]
  wire  io_in_writeResponse_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  io_in_writeResponse_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire  io_in_writeResponse_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  io_in_writeResponse_q_io_deq_valid; // @[Decoupled.scala 361:21]
  Queue_40 io_out_readAddress_q ( // @[Decoupled.scala 361:21]
    .clock(io_out_readAddress_q_clock),
    .reset(io_out_readAddress_q_reset),
    .io_enq_ready(io_out_readAddress_q_io_enq_ready),
    .io_enq_valid(io_out_readAddress_q_io_enq_valid),
    .io_enq_bits_addr(io_out_readAddress_q_io_enq_bits_addr),
    .io_enq_bits_len(io_out_readAddress_q_io_enq_bits_len),
    .io_enq_bits_cache(io_out_readAddress_q_io_enq_bits_cache),
    .io_deq_ready(io_out_readAddress_q_io_deq_ready),
    .io_deq_valid(io_out_readAddress_q_io_deq_valid),
    .io_deq_bits_id(io_out_readAddress_q_io_deq_bits_id),
    .io_deq_bits_addr(io_out_readAddress_q_io_deq_bits_addr),
    .io_deq_bits_len(io_out_readAddress_q_io_deq_bits_len),
    .io_deq_bits_size(io_out_readAddress_q_io_deq_bits_size),
    .io_deq_bits_burst(io_out_readAddress_q_io_deq_bits_burst),
    .io_deq_bits_lock(io_out_readAddress_q_io_deq_bits_lock),
    .io_deq_bits_cache(io_out_readAddress_q_io_deq_bits_cache),
    .io_deq_bits_prot(io_out_readAddress_q_io_deq_bits_prot),
    .io_deq_bits_qos(io_out_readAddress_q_io_deq_bits_qos)
  );
  Queue_40 io_out_writeAddress_q ( // @[Decoupled.scala 361:21]
    .clock(io_out_writeAddress_q_clock),
    .reset(io_out_writeAddress_q_reset),
    .io_enq_ready(io_out_writeAddress_q_io_enq_ready),
    .io_enq_valid(io_out_writeAddress_q_io_enq_valid),
    .io_enq_bits_addr(io_out_writeAddress_q_io_enq_bits_addr),
    .io_enq_bits_len(io_out_writeAddress_q_io_enq_bits_len),
    .io_enq_bits_cache(io_out_writeAddress_q_io_enq_bits_cache),
    .io_deq_ready(io_out_writeAddress_q_io_deq_ready),
    .io_deq_valid(io_out_writeAddress_q_io_deq_valid),
    .io_deq_bits_id(io_out_writeAddress_q_io_deq_bits_id),
    .io_deq_bits_addr(io_out_writeAddress_q_io_deq_bits_addr),
    .io_deq_bits_len(io_out_writeAddress_q_io_deq_bits_len),
    .io_deq_bits_size(io_out_writeAddress_q_io_deq_bits_size),
    .io_deq_bits_burst(io_out_writeAddress_q_io_deq_bits_burst),
    .io_deq_bits_lock(io_out_writeAddress_q_io_deq_bits_lock),
    .io_deq_bits_cache(io_out_writeAddress_q_io_deq_bits_cache),
    .io_deq_bits_prot(io_out_writeAddress_q_io_deq_bits_prot),
    .io_deq_bits_qos(io_out_writeAddress_q_io_deq_bits_qos)
  );
  Queue_42 io_out_writeData_q ( // @[Decoupled.scala 361:21]
    .clock(io_out_writeData_q_clock),
    .reset(io_out_writeData_q_reset),
    .io_enq_ready(io_out_writeData_q_io_enq_ready),
    .io_enq_valid(io_out_writeData_q_io_enq_valid),
    .io_enq_bits_data(io_out_writeData_q_io_enq_bits_data),
    .io_deq_ready(io_out_writeData_q_io_deq_ready),
    .io_deq_valid(io_out_writeData_q_io_deq_valid),
    .io_deq_bits_id(io_out_writeData_q_io_deq_bits_id),
    .io_deq_bits_data(io_out_writeData_q_io_deq_bits_data),
    .io_deq_bits_strb(io_out_writeData_q_io_deq_bits_strb)
  );
  Queue_38 io_in_readData_q ( // @[Decoupled.scala 361:21]
    .clock(io_in_readData_q_clock),
    .reset(io_in_readData_q_reset),
    .io_enq_ready(io_in_readData_q_io_enq_ready),
    .io_enq_valid(io_in_readData_q_io_enq_valid),
    .io_enq_bits_data(io_in_readData_q_io_enq_bits_data),
    .io_enq_bits_last(io_in_readData_q_io_enq_bits_last),
    .io_deq_ready(io_in_readData_q_io_deq_ready),
    .io_deq_valid(io_in_readData_q_io_deq_valid),
    .io_deq_bits_data(io_in_readData_q_io_deq_bits_data),
    .io_deq_bits_last(io_in_readData_q_io_deq_bits_last)
  );
  Queue_39 io_in_writeResponse_q ( // @[Decoupled.scala 361:21]
    .clock(io_in_writeResponse_q_clock),
    .reset(io_in_writeResponse_q_reset),
    .io_enq_ready(io_in_writeResponse_q_io_enq_ready),
    .io_enq_valid(io_in_writeResponse_q_io_enq_valid),
    .io_deq_ready(io_in_writeResponse_q_io_deq_ready),
    .io_deq_valid(io_in_writeResponse_q_io_deq_valid)
  );
  assign io_in_writeAddress_ready = io_out_writeAddress_q_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_in_writeData_ready = io_out_writeData_q_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_in_writeResponse_valid = io_in_writeResponse_q_io_deq_valid; // @[Queue.scala 18:23]
  assign io_in_readAddress_ready = io_out_readAddress_q_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_in_readData_valid = io_in_readData_q_io_deq_valid; // @[Queue.scala 17:18]
  assign io_in_readData_bits_data = io_in_readData_q_io_deq_bits_data; // @[Queue.scala 17:18]
  assign io_in_readData_bits_last = io_in_readData_q_io_deq_bits_last; // @[Queue.scala 17:18]
  assign io_out_writeAddress_valid = io_out_writeAddress_q_io_deq_valid; // @[Queue.scala 15:23]
  assign io_out_writeAddress_bits_id = io_out_writeAddress_q_io_deq_bits_id; // @[Queue.scala 15:23]
  assign io_out_writeAddress_bits_addr = io_out_writeAddress_q_io_deq_bits_addr; // @[Queue.scala 15:23]
  assign io_out_writeAddress_bits_len = io_out_writeAddress_q_io_deq_bits_len; // @[Queue.scala 15:23]
  assign io_out_writeAddress_bits_size = io_out_writeAddress_q_io_deq_bits_size; // @[Queue.scala 15:23]
  assign io_out_writeAddress_bits_burst = io_out_writeAddress_q_io_deq_bits_burst; // @[Queue.scala 15:23]
  assign io_out_writeAddress_bits_lock = io_out_writeAddress_q_io_deq_bits_lock; // @[Queue.scala 15:23]
  assign io_out_writeAddress_bits_cache = io_out_writeAddress_q_io_deq_bits_cache; // @[Queue.scala 15:23]
  assign io_out_writeAddress_bits_prot = io_out_writeAddress_q_io_deq_bits_prot; // @[Queue.scala 15:23]
  assign io_out_writeAddress_bits_qos = io_out_writeAddress_q_io_deq_bits_qos; // @[Queue.scala 15:23]
  assign io_out_writeData_valid = io_out_writeData_q_io_deq_valid; // @[Queue.scala 16:20]
  assign io_out_writeData_bits_id = io_out_writeData_q_io_deq_bits_id; // @[Queue.scala 16:20]
  assign io_out_writeData_bits_data = io_out_writeData_q_io_deq_bits_data; // @[Queue.scala 16:20]
  assign io_out_writeData_bits_strb = io_out_writeData_q_io_deq_bits_strb; // @[Queue.scala 16:20]
  assign io_out_writeResponse_ready = io_in_writeResponse_q_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_out_readAddress_valid = io_out_readAddress_q_io_deq_valid; // @[Queue.scala 14:22]
  assign io_out_readAddress_bits_id = io_out_readAddress_q_io_deq_bits_id; // @[Queue.scala 14:22]
  assign io_out_readAddress_bits_addr = io_out_readAddress_q_io_deq_bits_addr; // @[Queue.scala 14:22]
  assign io_out_readAddress_bits_len = io_out_readAddress_q_io_deq_bits_len; // @[Queue.scala 14:22]
  assign io_out_readAddress_bits_size = io_out_readAddress_q_io_deq_bits_size; // @[Queue.scala 14:22]
  assign io_out_readAddress_bits_burst = io_out_readAddress_q_io_deq_bits_burst; // @[Queue.scala 14:22]
  assign io_out_readAddress_bits_lock = io_out_readAddress_q_io_deq_bits_lock; // @[Queue.scala 14:22]
  assign io_out_readAddress_bits_cache = io_out_readAddress_q_io_deq_bits_cache; // @[Queue.scala 14:22]
  assign io_out_readAddress_bits_prot = io_out_readAddress_q_io_deq_bits_prot; // @[Queue.scala 14:22]
  assign io_out_readAddress_bits_qos = io_out_readAddress_q_io_deq_bits_qos; // @[Queue.scala 14:22]
  assign io_out_readData_ready = io_in_readData_q_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_out_readAddress_q_clock = clock;
  assign io_out_readAddress_q_reset = reset;
  assign io_out_readAddress_q_io_enq_valid = io_in_readAddress_valid; // @[Decoupled.scala 363:22]
  assign io_out_readAddress_q_io_enq_bits_addr = io_in_readAddress_bits_addr; // @[Decoupled.scala 364:21]
  assign io_out_readAddress_q_io_enq_bits_len = io_in_readAddress_bits_len; // @[Decoupled.scala 364:21]
  assign io_out_readAddress_q_io_enq_bits_cache = io_in_readAddress_bits_cache; // @[Decoupled.scala 364:21]
  assign io_out_readAddress_q_io_deq_ready = io_out_readAddress_ready; // @[Queue.scala 14:22]
  assign io_out_writeAddress_q_clock = clock;
  assign io_out_writeAddress_q_reset = reset;
  assign io_out_writeAddress_q_io_enq_valid = io_in_writeAddress_valid; // @[Decoupled.scala 363:22]
  assign io_out_writeAddress_q_io_enq_bits_addr = io_in_writeAddress_bits_addr; // @[Decoupled.scala 364:21]
  assign io_out_writeAddress_q_io_enq_bits_len = io_in_writeAddress_bits_len; // @[Decoupled.scala 364:21]
  assign io_out_writeAddress_q_io_enq_bits_cache = io_in_writeAddress_bits_cache; // @[Decoupled.scala 364:21]
  assign io_out_writeAddress_q_io_deq_ready = io_out_writeAddress_ready; // @[Queue.scala 15:23]
  assign io_out_writeData_q_clock = clock;
  assign io_out_writeData_q_reset = reset;
  assign io_out_writeData_q_io_enq_valid = io_in_writeData_valid; // @[Decoupled.scala 363:22]
  assign io_out_writeData_q_io_enq_bits_data = io_in_writeData_bits_data; // @[Decoupled.scala 364:21]
  assign io_out_writeData_q_io_deq_ready = io_out_writeData_ready; // @[Queue.scala 16:20]
  assign io_in_readData_q_clock = clock;
  assign io_in_readData_q_reset = reset;
  assign io_in_readData_q_io_enq_valid = io_out_readData_valid; // @[Decoupled.scala 363:22]
  assign io_in_readData_q_io_enq_bits_data = io_out_readData_bits_data; // @[Decoupled.scala 364:21]
  assign io_in_readData_q_io_enq_bits_last = io_out_readData_bits_last; // @[Decoupled.scala 364:21]
  assign io_in_readData_q_io_deq_ready = io_in_readData_ready; // @[Queue.scala 17:18]
  assign io_in_writeResponse_q_clock = clock;
  assign io_in_writeResponse_q_reset = reset;
  assign io_in_writeResponse_q_io_enq_valid = io_out_writeResponse_valid; // @[Decoupled.scala 363:22]
  assign io_in_writeResponse_q_io_deq_ready = io_in_writeResponse_ready; // @[Queue.scala 18:23]
endmodule
module AXIWrapperTCU(
  input          clock,
  input          reset,
  output         instruction_ready,
  input          instruction_valid,
  input  [3:0]   instruction_bits_opcode,
  input  [3:0]   instruction_bits_flags,
  input  [63:0]  instruction_bits_arguments,
  input          dram0_writeAddress_ready,
  output         dram0_writeAddress_valid,
  output [5:0]   dram0_writeAddress_bits_id,
  output [31:0]  dram0_writeAddress_bits_addr,
  output [7:0]   dram0_writeAddress_bits_len,
  output [2:0]   dram0_writeAddress_bits_size,
  output [1:0]   dram0_writeAddress_bits_burst,
  output [1:0]   dram0_writeAddress_bits_lock,
  output [3:0]   dram0_writeAddress_bits_cache,
  output [2:0]   dram0_writeAddress_bits_prot,
  output [3:0]   dram0_writeAddress_bits_qos,
  input          dram0_writeData_ready,
  output         dram0_writeData_valid,
  output [5:0]   dram0_writeData_bits_id,
  output [127:0] dram0_writeData_bits_data,
  output [15:0]  dram0_writeData_bits_strb,
  output         dram0_writeData_bits_last,
  output         dram0_writeResponse_ready,
  input          dram0_writeResponse_valid,
  input          dram0_readAddress_ready,
  output         dram0_readAddress_valid,
  output [5:0]   dram0_readAddress_bits_id,
  output [31:0]  dram0_readAddress_bits_addr,
  output [7:0]   dram0_readAddress_bits_len,
  output [2:0]   dram0_readAddress_bits_size,
  output [1:0]   dram0_readAddress_bits_burst,
  output [1:0]   dram0_readAddress_bits_lock,
  output [3:0]   dram0_readAddress_bits_cache,
  output [2:0]   dram0_readAddress_bits_prot,
  output [3:0]   dram0_readAddress_bits_qos,
  output         dram0_readData_ready,
  input          dram0_readData_valid,
  input  [127:0] dram0_readData_bits_data,
  input          dram1_writeAddress_ready,
  output         dram1_writeAddress_valid,
  output [5:0]   dram1_writeAddress_bits_id,
  output [31:0]  dram1_writeAddress_bits_addr,
  output [7:0]   dram1_writeAddress_bits_len,
  output [2:0]   dram1_writeAddress_bits_size,
  output [1:0]   dram1_writeAddress_bits_burst,
  output [1:0]   dram1_writeAddress_bits_lock,
  output [3:0]   dram1_writeAddress_bits_cache,
  output [2:0]   dram1_writeAddress_bits_prot,
  output [3:0]   dram1_writeAddress_bits_qos,
  input          dram1_writeData_ready,
  output         dram1_writeData_valid,
  output [5:0]   dram1_writeData_bits_id,
  output [127:0] dram1_writeData_bits_data,
  output [15:0]  dram1_writeData_bits_strb,
  output         dram1_writeData_bits_last,
  output         dram1_writeResponse_ready,
  input          dram1_writeResponse_valid,
  input          dram1_readAddress_ready,
  output         dram1_readAddress_valid,
  output [5:0]   dram1_readAddress_bits_id,
  output [31:0]  dram1_readAddress_bits_addr,
  output [7:0]   dram1_readAddress_bits_len,
  output [2:0]   dram1_readAddress_bits_size,
  output [1:0]   dram1_readAddress_bits_burst,
  output [1:0]   dram1_readAddress_bits_lock,
  output [3:0]   dram1_readAddress_bits_cache,
  output [2:0]   dram1_readAddress_bits_prot,
  output [3:0]   dram1_readAddress_bits_qos,
  output         dram1_readData_ready,
  input          dram1_readData_valid,
  input  [127:0] dram1_readData_bits_data
);
  wire  tcu_clock; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_reset; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_instruction_ready; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_instruction_valid; // @[AXIWrapperTCU.scala 32:19]
  wire [3:0] tcu_io_instruction_bits_opcode; // @[AXIWrapperTCU.scala 32:19]
  wire [3:0] tcu_io_instruction_bits_flags; // @[AXIWrapperTCU.scala 32:19]
  wire [63:0] tcu_io_instruction_bits_arguments; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram0_control_ready; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram0_control_valid; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram0_control_bits_write; // @[AXIWrapperTCU.scala 32:19]
  wire [20:0] tcu_io_dram0_control_bits_address; // @[AXIWrapperTCU.scala 32:19]
  wire [20:0] tcu_io_dram0_control_bits_size; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram0_dataIn_ready; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram0_dataIn_valid; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_0; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_1; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_2; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_3; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_4; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_5; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_6; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_7; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_8; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_9; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_10; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_11; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_12; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_13; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_14; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_15; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_16; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_17; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_18; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_19; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_20; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_21; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_22; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_23; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_24; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_25; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_26; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_27; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_28; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_29; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_30; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataIn_bits_31; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram0_dataOut_ready; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram0_dataOut_valid; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_0; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_1; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_2; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_3; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_4; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_5; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_6; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_7; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_8; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_9; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_10; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_11; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_12; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_13; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_14; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_15; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_16; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_17; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_18; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_19; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_20; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_21; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_22; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_23; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_24; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_25; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_26; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_27; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_28; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_29; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_30; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram0_dataOut_bits_31; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram1_control_ready; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram1_control_valid; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram1_control_bits_write; // @[AXIWrapperTCU.scala 32:19]
  wire [20:0] tcu_io_dram1_control_bits_address; // @[AXIWrapperTCU.scala 32:19]
  wire [20:0] tcu_io_dram1_control_bits_size; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram1_dataIn_ready; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram1_dataIn_valid; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_0; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_1; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_2; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_3; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_4; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_5; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_6; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_7; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_8; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_9; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_10; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_11; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_12; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_13; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_14; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_15; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_16; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_17; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_18; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_19; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_20; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_21; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_22; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_23; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_24; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_25; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_26; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_27; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_28; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_29; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_30; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataIn_bits_31; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram1_dataOut_ready; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_dram1_dataOut_valid; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_0; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_1; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_2; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_3; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_4; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_5; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_6; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_7; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_8; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_9; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_10; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_11; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_12; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_13; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_14; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_15; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_16; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_17; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_18; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_19; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_20; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_21; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_22; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_23; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_24; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_25; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_26; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_27; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_28; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_29; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_30; // @[AXIWrapperTCU.scala 32:19]
  wire [15:0] tcu_io_dram1_dataOut_bits_31; // @[AXIWrapperTCU.scala 32:19]
  wire [31:0] tcu_io_config_dram0AddressOffset; // @[AXIWrapperTCU.scala 32:19]
  wire [3:0] tcu_io_config_dram0CacheBehaviour; // @[AXIWrapperTCU.scala 32:19]
  wire [31:0] tcu_io_config_dram1AddressOffset; // @[AXIWrapperTCU.scala 32:19]
  wire [3:0] tcu_io_config_dram1CacheBehaviour; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_timeout; // @[AXIWrapperTCU.scala 32:19]
  wire  tcu_io_tracepoint; // @[AXIWrapperTCU.scala 32:19]
  wire [31:0] tcu_io_programCounter; // @[AXIWrapperTCU.scala 32:19]
  wire  dram0BoundarySplitter_clock; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_reset; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_writeAddress_ready; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_writeAddress_valid; // @[AXIWrapperTCU.scala 56:37]
  wire [5:0] dram0BoundarySplitter_io_in_writeAddress_bits_id; // @[AXIWrapperTCU.scala 56:37]
  wire [31:0] dram0BoundarySplitter_io_in_writeAddress_bits_addr; // @[AXIWrapperTCU.scala 56:37]
  wire [7:0] dram0BoundarySplitter_io_in_writeAddress_bits_len; // @[AXIWrapperTCU.scala 56:37]
  wire [2:0] dram0BoundarySplitter_io_in_writeAddress_bits_size; // @[AXIWrapperTCU.scala 56:37]
  wire [1:0] dram0BoundarySplitter_io_in_writeAddress_bits_burst; // @[AXIWrapperTCU.scala 56:37]
  wire [1:0] dram0BoundarySplitter_io_in_writeAddress_bits_lock; // @[AXIWrapperTCU.scala 56:37]
  wire [3:0] dram0BoundarySplitter_io_in_writeAddress_bits_cache; // @[AXIWrapperTCU.scala 56:37]
  wire [2:0] dram0BoundarySplitter_io_in_writeAddress_bits_prot; // @[AXIWrapperTCU.scala 56:37]
  wire [3:0] dram0BoundarySplitter_io_in_writeAddress_bits_qos; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_writeData_ready; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_writeData_valid; // @[AXIWrapperTCU.scala 56:37]
  wire [5:0] dram0BoundarySplitter_io_in_writeData_bits_id; // @[AXIWrapperTCU.scala 56:37]
  wire [127:0] dram0BoundarySplitter_io_in_writeData_bits_data; // @[AXIWrapperTCU.scala 56:37]
  wire [15:0] dram0BoundarySplitter_io_in_writeData_bits_strb; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_writeResponse_ready; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_writeResponse_valid; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_readAddress_ready; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_readAddress_valid; // @[AXIWrapperTCU.scala 56:37]
  wire [5:0] dram0BoundarySplitter_io_in_readAddress_bits_id; // @[AXIWrapperTCU.scala 56:37]
  wire [31:0] dram0BoundarySplitter_io_in_readAddress_bits_addr; // @[AXIWrapperTCU.scala 56:37]
  wire [7:0] dram0BoundarySplitter_io_in_readAddress_bits_len; // @[AXIWrapperTCU.scala 56:37]
  wire [2:0] dram0BoundarySplitter_io_in_readAddress_bits_size; // @[AXIWrapperTCU.scala 56:37]
  wire [1:0] dram0BoundarySplitter_io_in_readAddress_bits_burst; // @[AXIWrapperTCU.scala 56:37]
  wire [1:0] dram0BoundarySplitter_io_in_readAddress_bits_lock; // @[AXIWrapperTCU.scala 56:37]
  wire [3:0] dram0BoundarySplitter_io_in_readAddress_bits_cache; // @[AXIWrapperTCU.scala 56:37]
  wire [2:0] dram0BoundarySplitter_io_in_readAddress_bits_prot; // @[AXIWrapperTCU.scala 56:37]
  wire [3:0] dram0BoundarySplitter_io_in_readAddress_bits_qos; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_readData_ready; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_readData_valid; // @[AXIWrapperTCU.scala 56:37]
  wire [127:0] dram0BoundarySplitter_io_in_readData_bits_data; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_in_readData_bits_last; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_writeAddress_ready; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_writeAddress_valid; // @[AXIWrapperTCU.scala 56:37]
  wire [5:0] dram0BoundarySplitter_io_out_writeAddress_bits_id; // @[AXIWrapperTCU.scala 56:37]
  wire [31:0] dram0BoundarySplitter_io_out_writeAddress_bits_addr; // @[AXIWrapperTCU.scala 56:37]
  wire [7:0] dram0BoundarySplitter_io_out_writeAddress_bits_len; // @[AXIWrapperTCU.scala 56:37]
  wire [2:0] dram0BoundarySplitter_io_out_writeAddress_bits_size; // @[AXIWrapperTCU.scala 56:37]
  wire [1:0] dram0BoundarySplitter_io_out_writeAddress_bits_burst; // @[AXIWrapperTCU.scala 56:37]
  wire [1:0] dram0BoundarySplitter_io_out_writeAddress_bits_lock; // @[AXIWrapperTCU.scala 56:37]
  wire [3:0] dram0BoundarySplitter_io_out_writeAddress_bits_cache; // @[AXIWrapperTCU.scala 56:37]
  wire [2:0] dram0BoundarySplitter_io_out_writeAddress_bits_prot; // @[AXIWrapperTCU.scala 56:37]
  wire [3:0] dram0BoundarySplitter_io_out_writeAddress_bits_qos; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_writeData_ready; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_writeData_valid; // @[AXIWrapperTCU.scala 56:37]
  wire [5:0] dram0BoundarySplitter_io_out_writeData_bits_id; // @[AXIWrapperTCU.scala 56:37]
  wire [127:0] dram0BoundarySplitter_io_out_writeData_bits_data; // @[AXIWrapperTCU.scala 56:37]
  wire [15:0] dram0BoundarySplitter_io_out_writeData_bits_strb; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_writeData_bits_last; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_writeResponse_ready; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_writeResponse_valid; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_readAddress_ready; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_readAddress_valid; // @[AXIWrapperTCU.scala 56:37]
  wire [5:0] dram0BoundarySplitter_io_out_readAddress_bits_id; // @[AXIWrapperTCU.scala 56:37]
  wire [31:0] dram0BoundarySplitter_io_out_readAddress_bits_addr; // @[AXIWrapperTCU.scala 56:37]
  wire [7:0] dram0BoundarySplitter_io_out_readAddress_bits_len; // @[AXIWrapperTCU.scala 56:37]
  wire [2:0] dram0BoundarySplitter_io_out_readAddress_bits_size; // @[AXIWrapperTCU.scala 56:37]
  wire [1:0] dram0BoundarySplitter_io_out_readAddress_bits_burst; // @[AXIWrapperTCU.scala 56:37]
  wire [1:0] dram0BoundarySplitter_io_out_readAddress_bits_lock; // @[AXIWrapperTCU.scala 56:37]
  wire [3:0] dram0BoundarySplitter_io_out_readAddress_bits_cache; // @[AXIWrapperTCU.scala 56:37]
  wire [2:0] dram0BoundarySplitter_io_out_readAddress_bits_prot; // @[AXIWrapperTCU.scala 56:37]
  wire [3:0] dram0BoundarySplitter_io_out_readAddress_bits_qos; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_readData_ready; // @[AXIWrapperTCU.scala 56:37]
  wire  dram0BoundarySplitter_io_out_readData_valid; // @[AXIWrapperTCU.scala 56:37]
  wire [127:0] dram0BoundarySplitter_io_out_readData_bits_data; // @[AXIWrapperTCU.scala 56:37]
  wire  dram1BoundarySplitter_clock; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_reset; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_writeAddress_ready; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_writeAddress_valid; // @[AXIWrapperTCU.scala 60:37]
  wire [5:0] dram1BoundarySplitter_io_in_writeAddress_bits_id; // @[AXIWrapperTCU.scala 60:37]
  wire [31:0] dram1BoundarySplitter_io_in_writeAddress_bits_addr; // @[AXIWrapperTCU.scala 60:37]
  wire [7:0] dram1BoundarySplitter_io_in_writeAddress_bits_len; // @[AXIWrapperTCU.scala 60:37]
  wire [2:0] dram1BoundarySplitter_io_in_writeAddress_bits_size; // @[AXIWrapperTCU.scala 60:37]
  wire [1:0] dram1BoundarySplitter_io_in_writeAddress_bits_burst; // @[AXIWrapperTCU.scala 60:37]
  wire [1:0] dram1BoundarySplitter_io_in_writeAddress_bits_lock; // @[AXIWrapperTCU.scala 60:37]
  wire [3:0] dram1BoundarySplitter_io_in_writeAddress_bits_cache; // @[AXIWrapperTCU.scala 60:37]
  wire [2:0] dram1BoundarySplitter_io_in_writeAddress_bits_prot; // @[AXIWrapperTCU.scala 60:37]
  wire [3:0] dram1BoundarySplitter_io_in_writeAddress_bits_qos; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_writeData_ready; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_writeData_valid; // @[AXIWrapperTCU.scala 60:37]
  wire [5:0] dram1BoundarySplitter_io_in_writeData_bits_id; // @[AXIWrapperTCU.scala 60:37]
  wire [127:0] dram1BoundarySplitter_io_in_writeData_bits_data; // @[AXIWrapperTCU.scala 60:37]
  wire [15:0] dram1BoundarySplitter_io_in_writeData_bits_strb; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_writeResponse_ready; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_writeResponse_valid; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_readAddress_ready; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_readAddress_valid; // @[AXIWrapperTCU.scala 60:37]
  wire [5:0] dram1BoundarySplitter_io_in_readAddress_bits_id; // @[AXIWrapperTCU.scala 60:37]
  wire [31:0] dram1BoundarySplitter_io_in_readAddress_bits_addr; // @[AXIWrapperTCU.scala 60:37]
  wire [7:0] dram1BoundarySplitter_io_in_readAddress_bits_len; // @[AXIWrapperTCU.scala 60:37]
  wire [2:0] dram1BoundarySplitter_io_in_readAddress_bits_size; // @[AXIWrapperTCU.scala 60:37]
  wire [1:0] dram1BoundarySplitter_io_in_readAddress_bits_burst; // @[AXIWrapperTCU.scala 60:37]
  wire [1:0] dram1BoundarySplitter_io_in_readAddress_bits_lock; // @[AXIWrapperTCU.scala 60:37]
  wire [3:0] dram1BoundarySplitter_io_in_readAddress_bits_cache; // @[AXIWrapperTCU.scala 60:37]
  wire [2:0] dram1BoundarySplitter_io_in_readAddress_bits_prot; // @[AXIWrapperTCU.scala 60:37]
  wire [3:0] dram1BoundarySplitter_io_in_readAddress_bits_qos; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_readData_ready; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_readData_valid; // @[AXIWrapperTCU.scala 60:37]
  wire [127:0] dram1BoundarySplitter_io_in_readData_bits_data; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_in_readData_bits_last; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_writeAddress_ready; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_writeAddress_valid; // @[AXIWrapperTCU.scala 60:37]
  wire [5:0] dram1BoundarySplitter_io_out_writeAddress_bits_id; // @[AXIWrapperTCU.scala 60:37]
  wire [31:0] dram1BoundarySplitter_io_out_writeAddress_bits_addr; // @[AXIWrapperTCU.scala 60:37]
  wire [7:0] dram1BoundarySplitter_io_out_writeAddress_bits_len; // @[AXIWrapperTCU.scala 60:37]
  wire [2:0] dram1BoundarySplitter_io_out_writeAddress_bits_size; // @[AXIWrapperTCU.scala 60:37]
  wire [1:0] dram1BoundarySplitter_io_out_writeAddress_bits_burst; // @[AXIWrapperTCU.scala 60:37]
  wire [1:0] dram1BoundarySplitter_io_out_writeAddress_bits_lock; // @[AXIWrapperTCU.scala 60:37]
  wire [3:0] dram1BoundarySplitter_io_out_writeAddress_bits_cache; // @[AXIWrapperTCU.scala 60:37]
  wire [2:0] dram1BoundarySplitter_io_out_writeAddress_bits_prot; // @[AXIWrapperTCU.scala 60:37]
  wire [3:0] dram1BoundarySplitter_io_out_writeAddress_bits_qos; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_writeData_ready; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_writeData_valid; // @[AXIWrapperTCU.scala 60:37]
  wire [5:0] dram1BoundarySplitter_io_out_writeData_bits_id; // @[AXIWrapperTCU.scala 60:37]
  wire [127:0] dram1BoundarySplitter_io_out_writeData_bits_data; // @[AXIWrapperTCU.scala 60:37]
  wire [15:0] dram1BoundarySplitter_io_out_writeData_bits_strb; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_writeData_bits_last; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_writeResponse_ready; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_writeResponse_valid; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_readAddress_ready; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_readAddress_valid; // @[AXIWrapperTCU.scala 60:37]
  wire [5:0] dram1BoundarySplitter_io_out_readAddress_bits_id; // @[AXIWrapperTCU.scala 60:37]
  wire [31:0] dram1BoundarySplitter_io_out_readAddress_bits_addr; // @[AXIWrapperTCU.scala 60:37]
  wire [7:0] dram1BoundarySplitter_io_out_readAddress_bits_len; // @[AXIWrapperTCU.scala 60:37]
  wire [2:0] dram1BoundarySplitter_io_out_readAddress_bits_size; // @[AXIWrapperTCU.scala 60:37]
  wire [1:0] dram1BoundarySplitter_io_out_readAddress_bits_burst; // @[AXIWrapperTCU.scala 60:37]
  wire [1:0] dram1BoundarySplitter_io_out_readAddress_bits_lock; // @[AXIWrapperTCU.scala 60:37]
  wire [3:0] dram1BoundarySplitter_io_out_readAddress_bits_cache; // @[AXIWrapperTCU.scala 60:37]
  wire [2:0] dram1BoundarySplitter_io_out_readAddress_bits_prot; // @[AXIWrapperTCU.scala 60:37]
  wire [3:0] dram1BoundarySplitter_io_out_readAddress_bits_qos; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_readData_ready; // @[AXIWrapperTCU.scala 60:37]
  wire  dram1BoundarySplitter_io_out_readData_valid; // @[AXIWrapperTCU.scala 60:37]
  wire [127:0] dram1BoundarySplitter_io_out_readData_bits_data; // @[AXIWrapperTCU.scala 60:37]
  wire  dram0Converter_clock; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_reset; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_mem_control_ready; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_mem_control_valid; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_mem_control_bits_write; // @[AXIWrapperTCU.scala 65:30]
  wire [20:0] dram0Converter_io_mem_control_bits_address; // @[AXIWrapperTCU.scala 65:30]
  wire [20:0] dram0Converter_io_mem_control_bits_size; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_mem_dataIn_ready; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_mem_dataIn_valid; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_0; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_1; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_2; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_3; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_4; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_5; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_6; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_7; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_8; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_9; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_10; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_11; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_12; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_13; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_14; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_15; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_16; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_17; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_18; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_19; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_20; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_21; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_22; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_23; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_24; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_25; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_26; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_27; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_28; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_29; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_30; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataIn_bits_31; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_mem_dataOut_ready; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_mem_dataOut_valid; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_0; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_1; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_2; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_3; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_4; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_5; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_6; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_7; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_8; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_9; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_10; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_11; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_12; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_13; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_14; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_15; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_16; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_17; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_18; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_19; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_20; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_21; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_22; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_23; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_24; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_25; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_26; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_27; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_28; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_29; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_30; // @[AXIWrapperTCU.scala 65:30]
  wire [15:0] dram0Converter_io_mem_dataOut_bits_31; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_writeAddress_ready; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_writeAddress_valid; // @[AXIWrapperTCU.scala 65:30]
  wire [31:0] dram0Converter_io_axi_writeAddress_bits_addr; // @[AXIWrapperTCU.scala 65:30]
  wire [7:0] dram0Converter_io_axi_writeAddress_bits_len; // @[AXIWrapperTCU.scala 65:30]
  wire [3:0] dram0Converter_io_axi_writeAddress_bits_cache; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_writeData_ready; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_writeData_valid; // @[AXIWrapperTCU.scala 65:30]
  wire [127:0] dram0Converter_io_axi_writeData_bits_data; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_writeResponse_ready; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_writeResponse_valid; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_readAddress_ready; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_readAddress_valid; // @[AXIWrapperTCU.scala 65:30]
  wire [31:0] dram0Converter_io_axi_readAddress_bits_addr; // @[AXIWrapperTCU.scala 65:30]
  wire [7:0] dram0Converter_io_axi_readAddress_bits_len; // @[AXIWrapperTCU.scala 65:30]
  wire [3:0] dram0Converter_io_axi_readAddress_bits_cache; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_readData_ready; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_readData_valid; // @[AXIWrapperTCU.scala 65:30]
  wire [127:0] dram0Converter_io_axi_readData_bits_data; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_axi_readData_bits_last; // @[AXIWrapperTCU.scala 65:30]
  wire [31:0] dram0Converter_io_addressOffset; // @[AXIWrapperTCU.scala 65:30]
  wire [3:0] dram0Converter_io_cacheBehavior; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_timeout; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0Converter_io_tracepoint; // @[AXIWrapperTCU.scala 65:30]
  wire [31:0] dram0Converter_io_programCounter; // @[AXIWrapperTCU.scala 65:30]
  wire  dram0BoundarySplitter_io_in_q_clock; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_reset; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_writeAddress_ready; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_writeAddress_valid; // @[Queue.scala 23:19]
  wire [31:0] dram0BoundarySplitter_io_in_q_io_in_writeAddress_bits_addr; // @[Queue.scala 23:19]
  wire [7:0] dram0BoundarySplitter_io_in_q_io_in_writeAddress_bits_len; // @[Queue.scala 23:19]
  wire [3:0] dram0BoundarySplitter_io_in_q_io_in_writeAddress_bits_cache; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_writeData_ready; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_writeData_valid; // @[Queue.scala 23:19]
  wire [127:0] dram0BoundarySplitter_io_in_q_io_in_writeData_bits_data; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_writeResponse_ready; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_writeResponse_valid; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_readAddress_ready; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_readAddress_valid; // @[Queue.scala 23:19]
  wire [31:0] dram0BoundarySplitter_io_in_q_io_in_readAddress_bits_addr; // @[Queue.scala 23:19]
  wire [7:0] dram0BoundarySplitter_io_in_q_io_in_readAddress_bits_len; // @[Queue.scala 23:19]
  wire [3:0] dram0BoundarySplitter_io_in_q_io_in_readAddress_bits_cache; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_readData_ready; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_readData_valid; // @[Queue.scala 23:19]
  wire [127:0] dram0BoundarySplitter_io_in_q_io_in_readData_bits_data; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_in_readData_bits_last; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_writeAddress_ready; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_writeAddress_valid; // @[Queue.scala 23:19]
  wire [5:0] dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_id; // @[Queue.scala 23:19]
  wire [31:0] dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_addr; // @[Queue.scala 23:19]
  wire [7:0] dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_len; // @[Queue.scala 23:19]
  wire [2:0] dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_size; // @[Queue.scala 23:19]
  wire [1:0] dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_burst; // @[Queue.scala 23:19]
  wire [1:0] dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_lock; // @[Queue.scala 23:19]
  wire [3:0] dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_cache; // @[Queue.scala 23:19]
  wire [2:0] dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_prot; // @[Queue.scala 23:19]
  wire [3:0] dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_qos; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_writeData_ready; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_writeData_valid; // @[Queue.scala 23:19]
  wire [5:0] dram0BoundarySplitter_io_in_q_io_out_writeData_bits_id; // @[Queue.scala 23:19]
  wire [127:0] dram0BoundarySplitter_io_in_q_io_out_writeData_bits_data; // @[Queue.scala 23:19]
  wire [15:0] dram0BoundarySplitter_io_in_q_io_out_writeData_bits_strb; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_writeResponse_ready; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_writeResponse_valid; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_readAddress_ready; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_readAddress_valid; // @[Queue.scala 23:19]
  wire [5:0] dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_id; // @[Queue.scala 23:19]
  wire [31:0] dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_addr; // @[Queue.scala 23:19]
  wire [7:0] dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_len; // @[Queue.scala 23:19]
  wire [2:0] dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_size; // @[Queue.scala 23:19]
  wire [1:0] dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_burst; // @[Queue.scala 23:19]
  wire [1:0] dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_lock; // @[Queue.scala 23:19]
  wire [3:0] dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_cache; // @[Queue.scala 23:19]
  wire [2:0] dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_prot; // @[Queue.scala 23:19]
  wire [3:0] dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_qos; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_readData_ready; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_readData_valid; // @[Queue.scala 23:19]
  wire [127:0] dram0BoundarySplitter_io_in_q_io_out_readData_bits_data; // @[Queue.scala 23:19]
  wire  dram0BoundarySplitter_io_in_q_io_out_readData_bits_last; // @[Queue.scala 23:19]
  wire  dram1Converter_clock; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_reset; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_mem_control_ready; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_mem_control_valid; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_mem_control_bits_write; // @[AXIWrapperTCU.scala 82:30]
  wire [20:0] dram1Converter_io_mem_control_bits_address; // @[AXIWrapperTCU.scala 82:30]
  wire [20:0] dram1Converter_io_mem_control_bits_size; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_mem_dataIn_ready; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_mem_dataIn_valid; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_0; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_1; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_2; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_3; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_4; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_5; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_6; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_7; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_8; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_9; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_10; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_11; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_12; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_13; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_14; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_15; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_16; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_17; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_18; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_19; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_20; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_21; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_22; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_23; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_24; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_25; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_26; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_27; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_28; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_29; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_30; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataIn_bits_31; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_mem_dataOut_ready; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_mem_dataOut_valid; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_0; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_1; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_2; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_3; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_4; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_5; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_6; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_7; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_8; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_9; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_10; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_11; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_12; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_13; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_14; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_15; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_16; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_17; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_18; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_19; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_20; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_21; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_22; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_23; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_24; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_25; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_26; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_27; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_28; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_29; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_30; // @[AXIWrapperTCU.scala 82:30]
  wire [15:0] dram1Converter_io_mem_dataOut_bits_31; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_writeAddress_ready; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_writeAddress_valid; // @[AXIWrapperTCU.scala 82:30]
  wire [31:0] dram1Converter_io_axi_writeAddress_bits_addr; // @[AXIWrapperTCU.scala 82:30]
  wire [7:0] dram1Converter_io_axi_writeAddress_bits_len; // @[AXIWrapperTCU.scala 82:30]
  wire [3:0] dram1Converter_io_axi_writeAddress_bits_cache; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_writeData_ready; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_writeData_valid; // @[AXIWrapperTCU.scala 82:30]
  wire [127:0] dram1Converter_io_axi_writeData_bits_data; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_writeResponse_ready; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_writeResponse_valid; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_readAddress_ready; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_readAddress_valid; // @[AXIWrapperTCU.scala 82:30]
  wire [31:0] dram1Converter_io_axi_readAddress_bits_addr; // @[AXIWrapperTCU.scala 82:30]
  wire [7:0] dram1Converter_io_axi_readAddress_bits_len; // @[AXIWrapperTCU.scala 82:30]
  wire [3:0] dram1Converter_io_axi_readAddress_bits_cache; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_readData_ready; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_readData_valid; // @[AXIWrapperTCU.scala 82:30]
  wire [127:0] dram1Converter_io_axi_readData_bits_data; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_axi_readData_bits_last; // @[AXIWrapperTCU.scala 82:30]
  wire [31:0] dram1Converter_io_addressOffset; // @[AXIWrapperTCU.scala 82:30]
  wire [3:0] dram1Converter_io_cacheBehavior; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_timeout; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1Converter_io_tracepoint; // @[AXIWrapperTCU.scala 82:30]
  wire [31:0] dram1Converter_io_programCounter; // @[AXIWrapperTCU.scala 82:30]
  wire  dram1BoundarySplitter_io_in_q_clock; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_reset; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_writeAddress_ready; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_writeAddress_valid; // @[Queue.scala 23:19]
  wire [31:0] dram1BoundarySplitter_io_in_q_io_in_writeAddress_bits_addr; // @[Queue.scala 23:19]
  wire [7:0] dram1BoundarySplitter_io_in_q_io_in_writeAddress_bits_len; // @[Queue.scala 23:19]
  wire [3:0] dram1BoundarySplitter_io_in_q_io_in_writeAddress_bits_cache; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_writeData_ready; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_writeData_valid; // @[Queue.scala 23:19]
  wire [127:0] dram1BoundarySplitter_io_in_q_io_in_writeData_bits_data; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_writeResponse_ready; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_writeResponse_valid; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_readAddress_ready; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_readAddress_valid; // @[Queue.scala 23:19]
  wire [31:0] dram1BoundarySplitter_io_in_q_io_in_readAddress_bits_addr; // @[Queue.scala 23:19]
  wire [7:0] dram1BoundarySplitter_io_in_q_io_in_readAddress_bits_len; // @[Queue.scala 23:19]
  wire [3:0] dram1BoundarySplitter_io_in_q_io_in_readAddress_bits_cache; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_readData_ready; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_readData_valid; // @[Queue.scala 23:19]
  wire [127:0] dram1BoundarySplitter_io_in_q_io_in_readData_bits_data; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_in_readData_bits_last; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_writeAddress_ready; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_writeAddress_valid; // @[Queue.scala 23:19]
  wire [5:0] dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_id; // @[Queue.scala 23:19]
  wire [31:0] dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_addr; // @[Queue.scala 23:19]
  wire [7:0] dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_len; // @[Queue.scala 23:19]
  wire [2:0] dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_size; // @[Queue.scala 23:19]
  wire [1:0] dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_burst; // @[Queue.scala 23:19]
  wire [1:0] dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_lock; // @[Queue.scala 23:19]
  wire [3:0] dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_cache; // @[Queue.scala 23:19]
  wire [2:0] dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_prot; // @[Queue.scala 23:19]
  wire [3:0] dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_qos; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_writeData_ready; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_writeData_valid; // @[Queue.scala 23:19]
  wire [5:0] dram1BoundarySplitter_io_in_q_io_out_writeData_bits_id; // @[Queue.scala 23:19]
  wire [127:0] dram1BoundarySplitter_io_in_q_io_out_writeData_bits_data; // @[Queue.scala 23:19]
  wire [15:0] dram1BoundarySplitter_io_in_q_io_out_writeData_bits_strb; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_writeResponse_ready; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_writeResponse_valid; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_readAddress_ready; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_readAddress_valid; // @[Queue.scala 23:19]
  wire [5:0] dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_id; // @[Queue.scala 23:19]
  wire [31:0] dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_addr; // @[Queue.scala 23:19]
  wire [7:0] dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_len; // @[Queue.scala 23:19]
  wire [2:0] dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_size; // @[Queue.scala 23:19]
  wire [1:0] dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_burst; // @[Queue.scala 23:19]
  wire [1:0] dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_lock; // @[Queue.scala 23:19]
  wire [3:0] dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_cache; // @[Queue.scala 23:19]
  wire [2:0] dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_prot; // @[Queue.scala 23:19]
  wire [3:0] dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_qos; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_readData_ready; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_readData_valid; // @[Queue.scala 23:19]
  wire [127:0] dram1BoundarySplitter_io_in_q_io_out_readData_bits_data; // @[Queue.scala 23:19]
  wire  dram1BoundarySplitter_io_in_q_io_out_readData_bits_last; // @[Queue.scala 23:19]
  TCU tcu ( // @[AXIWrapperTCU.scala 32:19]
    .clock(tcu_clock),
    .reset(tcu_reset),
    .io_instruction_ready(tcu_io_instruction_ready),
    .io_instruction_valid(tcu_io_instruction_valid),
    .io_instruction_bits_opcode(tcu_io_instruction_bits_opcode),
    .io_instruction_bits_flags(tcu_io_instruction_bits_flags),
    .io_instruction_bits_arguments(tcu_io_instruction_bits_arguments),
    .io_dram0_control_ready(tcu_io_dram0_control_ready),
    .io_dram0_control_valid(tcu_io_dram0_control_valid),
    .io_dram0_control_bits_write(tcu_io_dram0_control_bits_write),
    .io_dram0_control_bits_address(tcu_io_dram0_control_bits_address),
    .io_dram0_control_bits_size(tcu_io_dram0_control_bits_size),
    .io_dram0_dataIn_ready(tcu_io_dram0_dataIn_ready),
    .io_dram0_dataIn_valid(tcu_io_dram0_dataIn_valid),
    .io_dram0_dataIn_bits_0(tcu_io_dram0_dataIn_bits_0),
    .io_dram0_dataIn_bits_1(tcu_io_dram0_dataIn_bits_1),
    .io_dram0_dataIn_bits_2(tcu_io_dram0_dataIn_bits_2),
    .io_dram0_dataIn_bits_3(tcu_io_dram0_dataIn_bits_3),
    .io_dram0_dataIn_bits_4(tcu_io_dram0_dataIn_bits_4),
    .io_dram0_dataIn_bits_5(tcu_io_dram0_dataIn_bits_5),
    .io_dram0_dataIn_bits_6(tcu_io_dram0_dataIn_bits_6),
    .io_dram0_dataIn_bits_7(tcu_io_dram0_dataIn_bits_7),
    .io_dram0_dataIn_bits_8(tcu_io_dram0_dataIn_bits_8),
    .io_dram0_dataIn_bits_9(tcu_io_dram0_dataIn_bits_9),
    .io_dram0_dataIn_bits_10(tcu_io_dram0_dataIn_bits_10),
    .io_dram0_dataIn_bits_11(tcu_io_dram0_dataIn_bits_11),
    .io_dram0_dataIn_bits_12(tcu_io_dram0_dataIn_bits_12),
    .io_dram0_dataIn_bits_13(tcu_io_dram0_dataIn_bits_13),
    .io_dram0_dataIn_bits_14(tcu_io_dram0_dataIn_bits_14),
    .io_dram0_dataIn_bits_15(tcu_io_dram0_dataIn_bits_15),
    .io_dram0_dataIn_bits_16(tcu_io_dram0_dataIn_bits_16),
    .io_dram0_dataIn_bits_17(tcu_io_dram0_dataIn_bits_17),
    .io_dram0_dataIn_bits_18(tcu_io_dram0_dataIn_bits_18),
    .io_dram0_dataIn_bits_19(tcu_io_dram0_dataIn_bits_19),
    .io_dram0_dataIn_bits_20(tcu_io_dram0_dataIn_bits_20),
    .io_dram0_dataIn_bits_21(tcu_io_dram0_dataIn_bits_21),
    .io_dram0_dataIn_bits_22(tcu_io_dram0_dataIn_bits_22),
    .io_dram0_dataIn_bits_23(tcu_io_dram0_dataIn_bits_23),
    .io_dram0_dataIn_bits_24(tcu_io_dram0_dataIn_bits_24),
    .io_dram0_dataIn_bits_25(tcu_io_dram0_dataIn_bits_25),
    .io_dram0_dataIn_bits_26(tcu_io_dram0_dataIn_bits_26),
    .io_dram0_dataIn_bits_27(tcu_io_dram0_dataIn_bits_27),
    .io_dram0_dataIn_bits_28(tcu_io_dram0_dataIn_bits_28),
    .io_dram0_dataIn_bits_29(tcu_io_dram0_dataIn_bits_29),
    .io_dram0_dataIn_bits_30(tcu_io_dram0_dataIn_bits_30),
    .io_dram0_dataIn_bits_31(tcu_io_dram0_dataIn_bits_31),
    .io_dram0_dataOut_ready(tcu_io_dram0_dataOut_ready),
    .io_dram0_dataOut_valid(tcu_io_dram0_dataOut_valid),
    .io_dram0_dataOut_bits_0(tcu_io_dram0_dataOut_bits_0),
    .io_dram0_dataOut_bits_1(tcu_io_dram0_dataOut_bits_1),
    .io_dram0_dataOut_bits_2(tcu_io_dram0_dataOut_bits_2),
    .io_dram0_dataOut_bits_3(tcu_io_dram0_dataOut_bits_3),
    .io_dram0_dataOut_bits_4(tcu_io_dram0_dataOut_bits_4),
    .io_dram0_dataOut_bits_5(tcu_io_dram0_dataOut_bits_5),
    .io_dram0_dataOut_bits_6(tcu_io_dram0_dataOut_bits_6),
    .io_dram0_dataOut_bits_7(tcu_io_dram0_dataOut_bits_7),
    .io_dram0_dataOut_bits_8(tcu_io_dram0_dataOut_bits_8),
    .io_dram0_dataOut_bits_9(tcu_io_dram0_dataOut_bits_9),
    .io_dram0_dataOut_bits_10(tcu_io_dram0_dataOut_bits_10),
    .io_dram0_dataOut_bits_11(tcu_io_dram0_dataOut_bits_11),
    .io_dram0_dataOut_bits_12(tcu_io_dram0_dataOut_bits_12),
    .io_dram0_dataOut_bits_13(tcu_io_dram0_dataOut_bits_13),
    .io_dram0_dataOut_bits_14(tcu_io_dram0_dataOut_bits_14),
    .io_dram0_dataOut_bits_15(tcu_io_dram0_dataOut_bits_15),
    .io_dram0_dataOut_bits_16(tcu_io_dram0_dataOut_bits_16),
    .io_dram0_dataOut_bits_17(tcu_io_dram0_dataOut_bits_17),
    .io_dram0_dataOut_bits_18(tcu_io_dram0_dataOut_bits_18),
    .io_dram0_dataOut_bits_19(tcu_io_dram0_dataOut_bits_19),
    .io_dram0_dataOut_bits_20(tcu_io_dram0_dataOut_bits_20),
    .io_dram0_dataOut_bits_21(tcu_io_dram0_dataOut_bits_21),
    .io_dram0_dataOut_bits_22(tcu_io_dram0_dataOut_bits_22),
    .io_dram0_dataOut_bits_23(tcu_io_dram0_dataOut_bits_23),
    .io_dram0_dataOut_bits_24(tcu_io_dram0_dataOut_bits_24),
    .io_dram0_dataOut_bits_25(tcu_io_dram0_dataOut_bits_25),
    .io_dram0_dataOut_bits_26(tcu_io_dram0_dataOut_bits_26),
    .io_dram0_dataOut_bits_27(tcu_io_dram0_dataOut_bits_27),
    .io_dram0_dataOut_bits_28(tcu_io_dram0_dataOut_bits_28),
    .io_dram0_dataOut_bits_29(tcu_io_dram0_dataOut_bits_29),
    .io_dram0_dataOut_bits_30(tcu_io_dram0_dataOut_bits_30),
    .io_dram0_dataOut_bits_31(tcu_io_dram0_dataOut_bits_31),
    .io_dram1_control_ready(tcu_io_dram1_control_ready),
    .io_dram1_control_valid(tcu_io_dram1_control_valid),
    .io_dram1_control_bits_write(tcu_io_dram1_control_bits_write),
    .io_dram1_control_bits_address(tcu_io_dram1_control_bits_address),
    .io_dram1_control_bits_size(tcu_io_dram1_control_bits_size),
    .io_dram1_dataIn_ready(tcu_io_dram1_dataIn_ready),
    .io_dram1_dataIn_valid(tcu_io_dram1_dataIn_valid),
    .io_dram1_dataIn_bits_0(tcu_io_dram1_dataIn_bits_0),
    .io_dram1_dataIn_bits_1(tcu_io_dram1_dataIn_bits_1),
    .io_dram1_dataIn_bits_2(tcu_io_dram1_dataIn_bits_2),
    .io_dram1_dataIn_bits_3(tcu_io_dram1_dataIn_bits_3),
    .io_dram1_dataIn_bits_4(tcu_io_dram1_dataIn_bits_4),
    .io_dram1_dataIn_bits_5(tcu_io_dram1_dataIn_bits_5),
    .io_dram1_dataIn_bits_6(tcu_io_dram1_dataIn_bits_6),
    .io_dram1_dataIn_bits_7(tcu_io_dram1_dataIn_bits_7),
    .io_dram1_dataIn_bits_8(tcu_io_dram1_dataIn_bits_8),
    .io_dram1_dataIn_bits_9(tcu_io_dram1_dataIn_bits_9),
    .io_dram1_dataIn_bits_10(tcu_io_dram1_dataIn_bits_10),
    .io_dram1_dataIn_bits_11(tcu_io_dram1_dataIn_bits_11),
    .io_dram1_dataIn_bits_12(tcu_io_dram1_dataIn_bits_12),
    .io_dram1_dataIn_bits_13(tcu_io_dram1_dataIn_bits_13),
    .io_dram1_dataIn_bits_14(tcu_io_dram1_dataIn_bits_14),
    .io_dram1_dataIn_bits_15(tcu_io_dram1_dataIn_bits_15),
    .io_dram1_dataIn_bits_16(tcu_io_dram1_dataIn_bits_16),
    .io_dram1_dataIn_bits_17(tcu_io_dram1_dataIn_bits_17),
    .io_dram1_dataIn_bits_18(tcu_io_dram1_dataIn_bits_18),
    .io_dram1_dataIn_bits_19(tcu_io_dram1_dataIn_bits_19),
    .io_dram1_dataIn_bits_20(tcu_io_dram1_dataIn_bits_20),
    .io_dram1_dataIn_bits_21(tcu_io_dram1_dataIn_bits_21),
    .io_dram1_dataIn_bits_22(tcu_io_dram1_dataIn_bits_22),
    .io_dram1_dataIn_bits_23(tcu_io_dram1_dataIn_bits_23),
    .io_dram1_dataIn_bits_24(tcu_io_dram1_dataIn_bits_24),
    .io_dram1_dataIn_bits_25(tcu_io_dram1_dataIn_bits_25),
    .io_dram1_dataIn_bits_26(tcu_io_dram1_dataIn_bits_26),
    .io_dram1_dataIn_bits_27(tcu_io_dram1_dataIn_bits_27),
    .io_dram1_dataIn_bits_28(tcu_io_dram1_dataIn_bits_28),
    .io_dram1_dataIn_bits_29(tcu_io_dram1_dataIn_bits_29),
    .io_dram1_dataIn_bits_30(tcu_io_dram1_dataIn_bits_30),
    .io_dram1_dataIn_bits_31(tcu_io_dram1_dataIn_bits_31),
    .io_dram1_dataOut_ready(tcu_io_dram1_dataOut_ready),
    .io_dram1_dataOut_valid(tcu_io_dram1_dataOut_valid),
    .io_dram1_dataOut_bits_0(tcu_io_dram1_dataOut_bits_0),
    .io_dram1_dataOut_bits_1(tcu_io_dram1_dataOut_bits_1),
    .io_dram1_dataOut_bits_2(tcu_io_dram1_dataOut_bits_2),
    .io_dram1_dataOut_bits_3(tcu_io_dram1_dataOut_bits_3),
    .io_dram1_dataOut_bits_4(tcu_io_dram1_dataOut_bits_4),
    .io_dram1_dataOut_bits_5(tcu_io_dram1_dataOut_bits_5),
    .io_dram1_dataOut_bits_6(tcu_io_dram1_dataOut_bits_6),
    .io_dram1_dataOut_bits_7(tcu_io_dram1_dataOut_bits_7),
    .io_dram1_dataOut_bits_8(tcu_io_dram1_dataOut_bits_8),
    .io_dram1_dataOut_bits_9(tcu_io_dram1_dataOut_bits_9),
    .io_dram1_dataOut_bits_10(tcu_io_dram1_dataOut_bits_10),
    .io_dram1_dataOut_bits_11(tcu_io_dram1_dataOut_bits_11),
    .io_dram1_dataOut_bits_12(tcu_io_dram1_dataOut_bits_12),
    .io_dram1_dataOut_bits_13(tcu_io_dram1_dataOut_bits_13),
    .io_dram1_dataOut_bits_14(tcu_io_dram1_dataOut_bits_14),
    .io_dram1_dataOut_bits_15(tcu_io_dram1_dataOut_bits_15),
    .io_dram1_dataOut_bits_16(tcu_io_dram1_dataOut_bits_16),
    .io_dram1_dataOut_bits_17(tcu_io_dram1_dataOut_bits_17),
    .io_dram1_dataOut_bits_18(tcu_io_dram1_dataOut_bits_18),
    .io_dram1_dataOut_bits_19(tcu_io_dram1_dataOut_bits_19),
    .io_dram1_dataOut_bits_20(tcu_io_dram1_dataOut_bits_20),
    .io_dram1_dataOut_bits_21(tcu_io_dram1_dataOut_bits_21),
    .io_dram1_dataOut_bits_22(tcu_io_dram1_dataOut_bits_22),
    .io_dram1_dataOut_bits_23(tcu_io_dram1_dataOut_bits_23),
    .io_dram1_dataOut_bits_24(tcu_io_dram1_dataOut_bits_24),
    .io_dram1_dataOut_bits_25(tcu_io_dram1_dataOut_bits_25),
    .io_dram1_dataOut_bits_26(tcu_io_dram1_dataOut_bits_26),
    .io_dram1_dataOut_bits_27(tcu_io_dram1_dataOut_bits_27),
    .io_dram1_dataOut_bits_28(tcu_io_dram1_dataOut_bits_28),
    .io_dram1_dataOut_bits_29(tcu_io_dram1_dataOut_bits_29),
    .io_dram1_dataOut_bits_30(tcu_io_dram1_dataOut_bits_30),
    .io_dram1_dataOut_bits_31(tcu_io_dram1_dataOut_bits_31),
    .io_config_dram0AddressOffset(tcu_io_config_dram0AddressOffset),
    .io_config_dram0CacheBehaviour(tcu_io_config_dram0CacheBehaviour),
    .io_config_dram1AddressOffset(tcu_io_config_dram1AddressOffset),
    .io_config_dram1CacheBehaviour(tcu_io_config_dram1CacheBehaviour),
    .io_timeout(tcu_io_timeout),
    .io_tracepoint(tcu_io_tracepoint),
    .io_programCounter(tcu_io_programCounter)
  );
  MemBoundarySplitter dram0BoundarySplitter ( // @[AXIWrapperTCU.scala 56:37]
    .clock(dram0BoundarySplitter_clock),
    .reset(dram0BoundarySplitter_reset),
    .io_in_writeAddress_ready(dram0BoundarySplitter_io_in_writeAddress_ready),
    .io_in_writeAddress_valid(dram0BoundarySplitter_io_in_writeAddress_valid),
    .io_in_writeAddress_bits_id(dram0BoundarySplitter_io_in_writeAddress_bits_id),
    .io_in_writeAddress_bits_addr(dram0BoundarySplitter_io_in_writeAddress_bits_addr),
    .io_in_writeAddress_bits_len(dram0BoundarySplitter_io_in_writeAddress_bits_len),
    .io_in_writeAddress_bits_size(dram0BoundarySplitter_io_in_writeAddress_bits_size),
    .io_in_writeAddress_bits_burst(dram0BoundarySplitter_io_in_writeAddress_bits_burst),
    .io_in_writeAddress_bits_lock(dram0BoundarySplitter_io_in_writeAddress_bits_lock),
    .io_in_writeAddress_bits_cache(dram0BoundarySplitter_io_in_writeAddress_bits_cache),
    .io_in_writeAddress_bits_prot(dram0BoundarySplitter_io_in_writeAddress_bits_prot),
    .io_in_writeAddress_bits_qos(dram0BoundarySplitter_io_in_writeAddress_bits_qos),
    .io_in_writeData_ready(dram0BoundarySplitter_io_in_writeData_ready),
    .io_in_writeData_valid(dram0BoundarySplitter_io_in_writeData_valid),
    .io_in_writeData_bits_id(dram0BoundarySplitter_io_in_writeData_bits_id),
    .io_in_writeData_bits_data(dram0BoundarySplitter_io_in_writeData_bits_data),
    .io_in_writeData_bits_strb(dram0BoundarySplitter_io_in_writeData_bits_strb),
    .io_in_writeResponse_ready(dram0BoundarySplitter_io_in_writeResponse_ready),
    .io_in_writeResponse_valid(dram0BoundarySplitter_io_in_writeResponse_valid),
    .io_in_readAddress_ready(dram0BoundarySplitter_io_in_readAddress_ready),
    .io_in_readAddress_valid(dram0BoundarySplitter_io_in_readAddress_valid),
    .io_in_readAddress_bits_id(dram0BoundarySplitter_io_in_readAddress_bits_id),
    .io_in_readAddress_bits_addr(dram0BoundarySplitter_io_in_readAddress_bits_addr),
    .io_in_readAddress_bits_len(dram0BoundarySplitter_io_in_readAddress_bits_len),
    .io_in_readAddress_bits_size(dram0BoundarySplitter_io_in_readAddress_bits_size),
    .io_in_readAddress_bits_burst(dram0BoundarySplitter_io_in_readAddress_bits_burst),
    .io_in_readAddress_bits_lock(dram0BoundarySplitter_io_in_readAddress_bits_lock),
    .io_in_readAddress_bits_cache(dram0BoundarySplitter_io_in_readAddress_bits_cache),
    .io_in_readAddress_bits_prot(dram0BoundarySplitter_io_in_readAddress_bits_prot),
    .io_in_readAddress_bits_qos(dram0BoundarySplitter_io_in_readAddress_bits_qos),
    .io_in_readData_ready(dram0BoundarySplitter_io_in_readData_ready),
    .io_in_readData_valid(dram0BoundarySplitter_io_in_readData_valid),
    .io_in_readData_bits_data(dram0BoundarySplitter_io_in_readData_bits_data),
    .io_in_readData_bits_last(dram0BoundarySplitter_io_in_readData_bits_last),
    .io_out_writeAddress_ready(dram0BoundarySplitter_io_out_writeAddress_ready),
    .io_out_writeAddress_valid(dram0BoundarySplitter_io_out_writeAddress_valid),
    .io_out_writeAddress_bits_id(dram0BoundarySplitter_io_out_writeAddress_bits_id),
    .io_out_writeAddress_bits_addr(dram0BoundarySplitter_io_out_writeAddress_bits_addr),
    .io_out_writeAddress_bits_len(dram0BoundarySplitter_io_out_writeAddress_bits_len),
    .io_out_writeAddress_bits_size(dram0BoundarySplitter_io_out_writeAddress_bits_size),
    .io_out_writeAddress_bits_burst(dram0BoundarySplitter_io_out_writeAddress_bits_burst),
    .io_out_writeAddress_bits_lock(dram0BoundarySplitter_io_out_writeAddress_bits_lock),
    .io_out_writeAddress_bits_cache(dram0BoundarySplitter_io_out_writeAddress_bits_cache),
    .io_out_writeAddress_bits_prot(dram0BoundarySplitter_io_out_writeAddress_bits_prot),
    .io_out_writeAddress_bits_qos(dram0BoundarySplitter_io_out_writeAddress_bits_qos),
    .io_out_writeData_ready(dram0BoundarySplitter_io_out_writeData_ready),
    .io_out_writeData_valid(dram0BoundarySplitter_io_out_writeData_valid),
    .io_out_writeData_bits_id(dram0BoundarySplitter_io_out_writeData_bits_id),
    .io_out_writeData_bits_data(dram0BoundarySplitter_io_out_writeData_bits_data),
    .io_out_writeData_bits_strb(dram0BoundarySplitter_io_out_writeData_bits_strb),
    .io_out_writeData_bits_last(dram0BoundarySplitter_io_out_writeData_bits_last),
    .io_out_writeResponse_ready(dram0BoundarySplitter_io_out_writeResponse_ready),
    .io_out_writeResponse_valid(dram0BoundarySplitter_io_out_writeResponse_valid),
    .io_out_readAddress_ready(dram0BoundarySplitter_io_out_readAddress_ready),
    .io_out_readAddress_valid(dram0BoundarySplitter_io_out_readAddress_valid),
    .io_out_readAddress_bits_id(dram0BoundarySplitter_io_out_readAddress_bits_id),
    .io_out_readAddress_bits_addr(dram0BoundarySplitter_io_out_readAddress_bits_addr),
    .io_out_readAddress_bits_len(dram0BoundarySplitter_io_out_readAddress_bits_len),
    .io_out_readAddress_bits_size(dram0BoundarySplitter_io_out_readAddress_bits_size),
    .io_out_readAddress_bits_burst(dram0BoundarySplitter_io_out_readAddress_bits_burst),
    .io_out_readAddress_bits_lock(dram0BoundarySplitter_io_out_readAddress_bits_lock),
    .io_out_readAddress_bits_cache(dram0BoundarySplitter_io_out_readAddress_bits_cache),
    .io_out_readAddress_bits_prot(dram0BoundarySplitter_io_out_readAddress_bits_prot),
    .io_out_readAddress_bits_qos(dram0BoundarySplitter_io_out_readAddress_bits_qos),
    .io_out_readData_ready(dram0BoundarySplitter_io_out_readData_ready),
    .io_out_readData_valid(dram0BoundarySplitter_io_out_readData_valid),
    .io_out_readData_bits_data(dram0BoundarySplitter_io_out_readData_bits_data)
  );
  MemBoundarySplitter dram1BoundarySplitter ( // @[AXIWrapperTCU.scala 60:37]
    .clock(dram1BoundarySplitter_clock),
    .reset(dram1BoundarySplitter_reset),
    .io_in_writeAddress_ready(dram1BoundarySplitter_io_in_writeAddress_ready),
    .io_in_writeAddress_valid(dram1BoundarySplitter_io_in_writeAddress_valid),
    .io_in_writeAddress_bits_id(dram1BoundarySplitter_io_in_writeAddress_bits_id),
    .io_in_writeAddress_bits_addr(dram1BoundarySplitter_io_in_writeAddress_bits_addr),
    .io_in_writeAddress_bits_len(dram1BoundarySplitter_io_in_writeAddress_bits_len),
    .io_in_writeAddress_bits_size(dram1BoundarySplitter_io_in_writeAddress_bits_size),
    .io_in_writeAddress_bits_burst(dram1BoundarySplitter_io_in_writeAddress_bits_burst),
    .io_in_writeAddress_bits_lock(dram1BoundarySplitter_io_in_writeAddress_bits_lock),
    .io_in_writeAddress_bits_cache(dram1BoundarySplitter_io_in_writeAddress_bits_cache),
    .io_in_writeAddress_bits_prot(dram1BoundarySplitter_io_in_writeAddress_bits_prot),
    .io_in_writeAddress_bits_qos(dram1BoundarySplitter_io_in_writeAddress_bits_qos),
    .io_in_writeData_ready(dram1BoundarySplitter_io_in_writeData_ready),
    .io_in_writeData_valid(dram1BoundarySplitter_io_in_writeData_valid),
    .io_in_writeData_bits_id(dram1BoundarySplitter_io_in_writeData_bits_id),
    .io_in_writeData_bits_data(dram1BoundarySplitter_io_in_writeData_bits_data),
    .io_in_writeData_bits_strb(dram1BoundarySplitter_io_in_writeData_bits_strb),
    .io_in_writeResponse_ready(dram1BoundarySplitter_io_in_writeResponse_ready),
    .io_in_writeResponse_valid(dram1BoundarySplitter_io_in_writeResponse_valid),
    .io_in_readAddress_ready(dram1BoundarySplitter_io_in_readAddress_ready),
    .io_in_readAddress_valid(dram1BoundarySplitter_io_in_readAddress_valid),
    .io_in_readAddress_bits_id(dram1BoundarySplitter_io_in_readAddress_bits_id),
    .io_in_readAddress_bits_addr(dram1BoundarySplitter_io_in_readAddress_bits_addr),
    .io_in_readAddress_bits_len(dram1BoundarySplitter_io_in_readAddress_bits_len),
    .io_in_readAddress_bits_size(dram1BoundarySplitter_io_in_readAddress_bits_size),
    .io_in_readAddress_bits_burst(dram1BoundarySplitter_io_in_readAddress_bits_burst),
    .io_in_readAddress_bits_lock(dram1BoundarySplitter_io_in_readAddress_bits_lock),
    .io_in_readAddress_bits_cache(dram1BoundarySplitter_io_in_readAddress_bits_cache),
    .io_in_readAddress_bits_prot(dram1BoundarySplitter_io_in_readAddress_bits_prot),
    .io_in_readAddress_bits_qos(dram1BoundarySplitter_io_in_readAddress_bits_qos),
    .io_in_readData_ready(dram1BoundarySplitter_io_in_readData_ready),
    .io_in_readData_valid(dram1BoundarySplitter_io_in_readData_valid),
    .io_in_readData_bits_data(dram1BoundarySplitter_io_in_readData_bits_data),
    .io_in_readData_bits_last(dram1BoundarySplitter_io_in_readData_bits_last),
    .io_out_writeAddress_ready(dram1BoundarySplitter_io_out_writeAddress_ready),
    .io_out_writeAddress_valid(dram1BoundarySplitter_io_out_writeAddress_valid),
    .io_out_writeAddress_bits_id(dram1BoundarySplitter_io_out_writeAddress_bits_id),
    .io_out_writeAddress_bits_addr(dram1BoundarySplitter_io_out_writeAddress_bits_addr),
    .io_out_writeAddress_bits_len(dram1BoundarySplitter_io_out_writeAddress_bits_len),
    .io_out_writeAddress_bits_size(dram1BoundarySplitter_io_out_writeAddress_bits_size),
    .io_out_writeAddress_bits_burst(dram1BoundarySplitter_io_out_writeAddress_bits_burst),
    .io_out_writeAddress_bits_lock(dram1BoundarySplitter_io_out_writeAddress_bits_lock),
    .io_out_writeAddress_bits_cache(dram1BoundarySplitter_io_out_writeAddress_bits_cache),
    .io_out_writeAddress_bits_prot(dram1BoundarySplitter_io_out_writeAddress_bits_prot),
    .io_out_writeAddress_bits_qos(dram1BoundarySplitter_io_out_writeAddress_bits_qos),
    .io_out_writeData_ready(dram1BoundarySplitter_io_out_writeData_ready),
    .io_out_writeData_valid(dram1BoundarySplitter_io_out_writeData_valid),
    .io_out_writeData_bits_id(dram1BoundarySplitter_io_out_writeData_bits_id),
    .io_out_writeData_bits_data(dram1BoundarySplitter_io_out_writeData_bits_data),
    .io_out_writeData_bits_strb(dram1BoundarySplitter_io_out_writeData_bits_strb),
    .io_out_writeData_bits_last(dram1BoundarySplitter_io_out_writeData_bits_last),
    .io_out_writeResponse_ready(dram1BoundarySplitter_io_out_writeResponse_ready),
    .io_out_writeResponse_valid(dram1BoundarySplitter_io_out_writeResponse_valid),
    .io_out_readAddress_ready(dram1BoundarySplitter_io_out_readAddress_ready),
    .io_out_readAddress_valid(dram1BoundarySplitter_io_out_readAddress_valid),
    .io_out_readAddress_bits_id(dram1BoundarySplitter_io_out_readAddress_bits_id),
    .io_out_readAddress_bits_addr(dram1BoundarySplitter_io_out_readAddress_bits_addr),
    .io_out_readAddress_bits_len(dram1BoundarySplitter_io_out_readAddress_bits_len),
    .io_out_readAddress_bits_size(dram1BoundarySplitter_io_out_readAddress_bits_size),
    .io_out_readAddress_bits_burst(dram1BoundarySplitter_io_out_readAddress_bits_burst),
    .io_out_readAddress_bits_lock(dram1BoundarySplitter_io_out_readAddress_bits_lock),
    .io_out_readAddress_bits_cache(dram1BoundarySplitter_io_out_readAddress_bits_cache),
    .io_out_readAddress_bits_prot(dram1BoundarySplitter_io_out_readAddress_bits_prot),
    .io_out_readAddress_bits_qos(dram1BoundarySplitter_io_out_readAddress_bits_qos),
    .io_out_readData_ready(dram1BoundarySplitter_io_out_readData_ready),
    .io_out_readData_valid(dram1BoundarySplitter_io_out_readData_valid),
    .io_out_readData_bits_data(dram1BoundarySplitter_io_out_readData_bits_data)
  );
  Converter dram0Converter ( // @[AXIWrapperTCU.scala 65:30]
    .clock(dram0Converter_clock),
    .reset(dram0Converter_reset),
    .io_mem_control_ready(dram0Converter_io_mem_control_ready),
    .io_mem_control_valid(dram0Converter_io_mem_control_valid),
    .io_mem_control_bits_write(dram0Converter_io_mem_control_bits_write),
    .io_mem_control_bits_address(dram0Converter_io_mem_control_bits_address),
    .io_mem_control_bits_size(dram0Converter_io_mem_control_bits_size),
    .io_mem_dataIn_ready(dram0Converter_io_mem_dataIn_ready),
    .io_mem_dataIn_valid(dram0Converter_io_mem_dataIn_valid),
    .io_mem_dataIn_bits_0(dram0Converter_io_mem_dataIn_bits_0),
    .io_mem_dataIn_bits_1(dram0Converter_io_mem_dataIn_bits_1),
    .io_mem_dataIn_bits_2(dram0Converter_io_mem_dataIn_bits_2),
    .io_mem_dataIn_bits_3(dram0Converter_io_mem_dataIn_bits_3),
    .io_mem_dataIn_bits_4(dram0Converter_io_mem_dataIn_bits_4),
    .io_mem_dataIn_bits_5(dram0Converter_io_mem_dataIn_bits_5),
    .io_mem_dataIn_bits_6(dram0Converter_io_mem_dataIn_bits_6),
    .io_mem_dataIn_bits_7(dram0Converter_io_mem_dataIn_bits_7),
    .io_mem_dataIn_bits_8(dram0Converter_io_mem_dataIn_bits_8),
    .io_mem_dataIn_bits_9(dram0Converter_io_mem_dataIn_bits_9),
    .io_mem_dataIn_bits_10(dram0Converter_io_mem_dataIn_bits_10),
    .io_mem_dataIn_bits_11(dram0Converter_io_mem_dataIn_bits_11),
    .io_mem_dataIn_bits_12(dram0Converter_io_mem_dataIn_bits_12),
    .io_mem_dataIn_bits_13(dram0Converter_io_mem_dataIn_bits_13),
    .io_mem_dataIn_bits_14(dram0Converter_io_mem_dataIn_bits_14),
    .io_mem_dataIn_bits_15(dram0Converter_io_mem_dataIn_bits_15),
    .io_mem_dataIn_bits_16(dram0Converter_io_mem_dataIn_bits_16),
    .io_mem_dataIn_bits_17(dram0Converter_io_mem_dataIn_bits_17),
    .io_mem_dataIn_bits_18(dram0Converter_io_mem_dataIn_bits_18),
    .io_mem_dataIn_bits_19(dram0Converter_io_mem_dataIn_bits_19),
    .io_mem_dataIn_bits_20(dram0Converter_io_mem_dataIn_bits_20),
    .io_mem_dataIn_bits_21(dram0Converter_io_mem_dataIn_bits_21),
    .io_mem_dataIn_bits_22(dram0Converter_io_mem_dataIn_bits_22),
    .io_mem_dataIn_bits_23(dram0Converter_io_mem_dataIn_bits_23),
    .io_mem_dataIn_bits_24(dram0Converter_io_mem_dataIn_bits_24),
    .io_mem_dataIn_bits_25(dram0Converter_io_mem_dataIn_bits_25),
    .io_mem_dataIn_bits_26(dram0Converter_io_mem_dataIn_bits_26),
    .io_mem_dataIn_bits_27(dram0Converter_io_mem_dataIn_bits_27),
    .io_mem_dataIn_bits_28(dram0Converter_io_mem_dataIn_bits_28),
    .io_mem_dataIn_bits_29(dram0Converter_io_mem_dataIn_bits_29),
    .io_mem_dataIn_bits_30(dram0Converter_io_mem_dataIn_bits_30),
    .io_mem_dataIn_bits_31(dram0Converter_io_mem_dataIn_bits_31),
    .io_mem_dataOut_ready(dram0Converter_io_mem_dataOut_ready),
    .io_mem_dataOut_valid(dram0Converter_io_mem_dataOut_valid),
    .io_mem_dataOut_bits_0(dram0Converter_io_mem_dataOut_bits_0),
    .io_mem_dataOut_bits_1(dram0Converter_io_mem_dataOut_bits_1),
    .io_mem_dataOut_bits_2(dram0Converter_io_mem_dataOut_bits_2),
    .io_mem_dataOut_bits_3(dram0Converter_io_mem_dataOut_bits_3),
    .io_mem_dataOut_bits_4(dram0Converter_io_mem_dataOut_bits_4),
    .io_mem_dataOut_bits_5(dram0Converter_io_mem_dataOut_bits_5),
    .io_mem_dataOut_bits_6(dram0Converter_io_mem_dataOut_bits_6),
    .io_mem_dataOut_bits_7(dram0Converter_io_mem_dataOut_bits_7),
    .io_mem_dataOut_bits_8(dram0Converter_io_mem_dataOut_bits_8),
    .io_mem_dataOut_bits_9(dram0Converter_io_mem_dataOut_bits_9),
    .io_mem_dataOut_bits_10(dram0Converter_io_mem_dataOut_bits_10),
    .io_mem_dataOut_bits_11(dram0Converter_io_mem_dataOut_bits_11),
    .io_mem_dataOut_bits_12(dram0Converter_io_mem_dataOut_bits_12),
    .io_mem_dataOut_bits_13(dram0Converter_io_mem_dataOut_bits_13),
    .io_mem_dataOut_bits_14(dram0Converter_io_mem_dataOut_bits_14),
    .io_mem_dataOut_bits_15(dram0Converter_io_mem_dataOut_bits_15),
    .io_mem_dataOut_bits_16(dram0Converter_io_mem_dataOut_bits_16),
    .io_mem_dataOut_bits_17(dram0Converter_io_mem_dataOut_bits_17),
    .io_mem_dataOut_bits_18(dram0Converter_io_mem_dataOut_bits_18),
    .io_mem_dataOut_bits_19(dram0Converter_io_mem_dataOut_bits_19),
    .io_mem_dataOut_bits_20(dram0Converter_io_mem_dataOut_bits_20),
    .io_mem_dataOut_bits_21(dram0Converter_io_mem_dataOut_bits_21),
    .io_mem_dataOut_bits_22(dram0Converter_io_mem_dataOut_bits_22),
    .io_mem_dataOut_bits_23(dram0Converter_io_mem_dataOut_bits_23),
    .io_mem_dataOut_bits_24(dram0Converter_io_mem_dataOut_bits_24),
    .io_mem_dataOut_bits_25(dram0Converter_io_mem_dataOut_bits_25),
    .io_mem_dataOut_bits_26(dram0Converter_io_mem_dataOut_bits_26),
    .io_mem_dataOut_bits_27(dram0Converter_io_mem_dataOut_bits_27),
    .io_mem_dataOut_bits_28(dram0Converter_io_mem_dataOut_bits_28),
    .io_mem_dataOut_bits_29(dram0Converter_io_mem_dataOut_bits_29),
    .io_mem_dataOut_bits_30(dram0Converter_io_mem_dataOut_bits_30),
    .io_mem_dataOut_bits_31(dram0Converter_io_mem_dataOut_bits_31),
    .io_axi_writeAddress_ready(dram0Converter_io_axi_writeAddress_ready),
    .io_axi_writeAddress_valid(dram0Converter_io_axi_writeAddress_valid),
    .io_axi_writeAddress_bits_addr(dram0Converter_io_axi_writeAddress_bits_addr),
    .io_axi_writeAddress_bits_len(dram0Converter_io_axi_writeAddress_bits_len),
    .io_axi_writeAddress_bits_cache(dram0Converter_io_axi_writeAddress_bits_cache),
    .io_axi_writeData_ready(dram0Converter_io_axi_writeData_ready),
    .io_axi_writeData_valid(dram0Converter_io_axi_writeData_valid),
    .io_axi_writeData_bits_data(dram0Converter_io_axi_writeData_bits_data),
    .io_axi_writeResponse_ready(dram0Converter_io_axi_writeResponse_ready),
    .io_axi_writeResponse_valid(dram0Converter_io_axi_writeResponse_valid),
    .io_axi_readAddress_ready(dram0Converter_io_axi_readAddress_ready),
    .io_axi_readAddress_valid(dram0Converter_io_axi_readAddress_valid),
    .io_axi_readAddress_bits_addr(dram0Converter_io_axi_readAddress_bits_addr),
    .io_axi_readAddress_bits_len(dram0Converter_io_axi_readAddress_bits_len),
    .io_axi_readAddress_bits_cache(dram0Converter_io_axi_readAddress_bits_cache),
    .io_axi_readData_ready(dram0Converter_io_axi_readData_ready),
    .io_axi_readData_valid(dram0Converter_io_axi_readData_valid),
    .io_axi_readData_bits_data(dram0Converter_io_axi_readData_bits_data),
    .io_axi_readData_bits_last(dram0Converter_io_axi_readData_bits_last),
    .io_addressOffset(dram0Converter_io_addressOffset),
    .io_cacheBehavior(dram0Converter_io_cacheBehavior),
    .io_timeout(dram0Converter_io_timeout),
    .io_tracepoint(dram0Converter_io_tracepoint),
    .io_programCounter(dram0Converter_io_programCounter)
  );
  Queue_45 dram0BoundarySplitter_io_in_q ( // @[Queue.scala 23:19]
    .clock(dram0BoundarySplitter_io_in_q_clock),
    .reset(dram0BoundarySplitter_io_in_q_reset),
    .io_in_writeAddress_ready(dram0BoundarySplitter_io_in_q_io_in_writeAddress_ready),
    .io_in_writeAddress_valid(dram0BoundarySplitter_io_in_q_io_in_writeAddress_valid),
    .io_in_writeAddress_bits_addr(dram0BoundarySplitter_io_in_q_io_in_writeAddress_bits_addr),
    .io_in_writeAddress_bits_len(dram0BoundarySplitter_io_in_q_io_in_writeAddress_bits_len),
    .io_in_writeAddress_bits_cache(dram0BoundarySplitter_io_in_q_io_in_writeAddress_bits_cache),
    .io_in_writeData_ready(dram0BoundarySplitter_io_in_q_io_in_writeData_ready),
    .io_in_writeData_valid(dram0BoundarySplitter_io_in_q_io_in_writeData_valid),
    .io_in_writeData_bits_data(dram0BoundarySplitter_io_in_q_io_in_writeData_bits_data),
    .io_in_writeResponse_ready(dram0BoundarySplitter_io_in_q_io_in_writeResponse_ready),
    .io_in_writeResponse_valid(dram0BoundarySplitter_io_in_q_io_in_writeResponse_valid),
    .io_in_readAddress_ready(dram0BoundarySplitter_io_in_q_io_in_readAddress_ready),
    .io_in_readAddress_valid(dram0BoundarySplitter_io_in_q_io_in_readAddress_valid),
    .io_in_readAddress_bits_addr(dram0BoundarySplitter_io_in_q_io_in_readAddress_bits_addr),
    .io_in_readAddress_bits_len(dram0BoundarySplitter_io_in_q_io_in_readAddress_bits_len),
    .io_in_readAddress_bits_cache(dram0BoundarySplitter_io_in_q_io_in_readAddress_bits_cache),
    .io_in_readData_ready(dram0BoundarySplitter_io_in_q_io_in_readData_ready),
    .io_in_readData_valid(dram0BoundarySplitter_io_in_q_io_in_readData_valid),
    .io_in_readData_bits_data(dram0BoundarySplitter_io_in_q_io_in_readData_bits_data),
    .io_in_readData_bits_last(dram0BoundarySplitter_io_in_q_io_in_readData_bits_last),
    .io_out_writeAddress_ready(dram0BoundarySplitter_io_in_q_io_out_writeAddress_ready),
    .io_out_writeAddress_valid(dram0BoundarySplitter_io_in_q_io_out_writeAddress_valid),
    .io_out_writeAddress_bits_id(dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_id),
    .io_out_writeAddress_bits_addr(dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_addr),
    .io_out_writeAddress_bits_len(dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_len),
    .io_out_writeAddress_bits_size(dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_size),
    .io_out_writeAddress_bits_burst(dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_burst),
    .io_out_writeAddress_bits_lock(dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_lock),
    .io_out_writeAddress_bits_cache(dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_cache),
    .io_out_writeAddress_bits_prot(dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_prot),
    .io_out_writeAddress_bits_qos(dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_qos),
    .io_out_writeData_ready(dram0BoundarySplitter_io_in_q_io_out_writeData_ready),
    .io_out_writeData_valid(dram0BoundarySplitter_io_in_q_io_out_writeData_valid),
    .io_out_writeData_bits_id(dram0BoundarySplitter_io_in_q_io_out_writeData_bits_id),
    .io_out_writeData_bits_data(dram0BoundarySplitter_io_in_q_io_out_writeData_bits_data),
    .io_out_writeData_bits_strb(dram0BoundarySplitter_io_in_q_io_out_writeData_bits_strb),
    .io_out_writeResponse_ready(dram0BoundarySplitter_io_in_q_io_out_writeResponse_ready),
    .io_out_writeResponse_valid(dram0BoundarySplitter_io_in_q_io_out_writeResponse_valid),
    .io_out_readAddress_ready(dram0BoundarySplitter_io_in_q_io_out_readAddress_ready),
    .io_out_readAddress_valid(dram0BoundarySplitter_io_in_q_io_out_readAddress_valid),
    .io_out_readAddress_bits_id(dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_id),
    .io_out_readAddress_bits_addr(dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_addr),
    .io_out_readAddress_bits_len(dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_len),
    .io_out_readAddress_bits_size(dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_size),
    .io_out_readAddress_bits_burst(dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_burst),
    .io_out_readAddress_bits_lock(dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_lock),
    .io_out_readAddress_bits_cache(dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_cache),
    .io_out_readAddress_bits_prot(dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_prot),
    .io_out_readAddress_bits_qos(dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_qos),
    .io_out_readData_ready(dram0BoundarySplitter_io_in_q_io_out_readData_ready),
    .io_out_readData_valid(dram0BoundarySplitter_io_in_q_io_out_readData_valid),
    .io_out_readData_bits_data(dram0BoundarySplitter_io_in_q_io_out_readData_bits_data),
    .io_out_readData_bits_last(dram0BoundarySplitter_io_in_q_io_out_readData_bits_last)
  );
  Converter dram1Converter ( // @[AXIWrapperTCU.scala 82:30]
    .clock(dram1Converter_clock),
    .reset(dram1Converter_reset),
    .io_mem_control_ready(dram1Converter_io_mem_control_ready),
    .io_mem_control_valid(dram1Converter_io_mem_control_valid),
    .io_mem_control_bits_write(dram1Converter_io_mem_control_bits_write),
    .io_mem_control_bits_address(dram1Converter_io_mem_control_bits_address),
    .io_mem_control_bits_size(dram1Converter_io_mem_control_bits_size),
    .io_mem_dataIn_ready(dram1Converter_io_mem_dataIn_ready),
    .io_mem_dataIn_valid(dram1Converter_io_mem_dataIn_valid),
    .io_mem_dataIn_bits_0(dram1Converter_io_mem_dataIn_bits_0),
    .io_mem_dataIn_bits_1(dram1Converter_io_mem_dataIn_bits_1),
    .io_mem_dataIn_bits_2(dram1Converter_io_mem_dataIn_bits_2),
    .io_mem_dataIn_bits_3(dram1Converter_io_mem_dataIn_bits_3),
    .io_mem_dataIn_bits_4(dram1Converter_io_mem_dataIn_bits_4),
    .io_mem_dataIn_bits_5(dram1Converter_io_mem_dataIn_bits_5),
    .io_mem_dataIn_bits_6(dram1Converter_io_mem_dataIn_bits_6),
    .io_mem_dataIn_bits_7(dram1Converter_io_mem_dataIn_bits_7),
    .io_mem_dataIn_bits_8(dram1Converter_io_mem_dataIn_bits_8),
    .io_mem_dataIn_bits_9(dram1Converter_io_mem_dataIn_bits_9),
    .io_mem_dataIn_bits_10(dram1Converter_io_mem_dataIn_bits_10),
    .io_mem_dataIn_bits_11(dram1Converter_io_mem_dataIn_bits_11),
    .io_mem_dataIn_bits_12(dram1Converter_io_mem_dataIn_bits_12),
    .io_mem_dataIn_bits_13(dram1Converter_io_mem_dataIn_bits_13),
    .io_mem_dataIn_bits_14(dram1Converter_io_mem_dataIn_bits_14),
    .io_mem_dataIn_bits_15(dram1Converter_io_mem_dataIn_bits_15),
    .io_mem_dataIn_bits_16(dram1Converter_io_mem_dataIn_bits_16),
    .io_mem_dataIn_bits_17(dram1Converter_io_mem_dataIn_bits_17),
    .io_mem_dataIn_bits_18(dram1Converter_io_mem_dataIn_bits_18),
    .io_mem_dataIn_bits_19(dram1Converter_io_mem_dataIn_bits_19),
    .io_mem_dataIn_bits_20(dram1Converter_io_mem_dataIn_bits_20),
    .io_mem_dataIn_bits_21(dram1Converter_io_mem_dataIn_bits_21),
    .io_mem_dataIn_bits_22(dram1Converter_io_mem_dataIn_bits_22),
    .io_mem_dataIn_bits_23(dram1Converter_io_mem_dataIn_bits_23),
    .io_mem_dataIn_bits_24(dram1Converter_io_mem_dataIn_bits_24),
    .io_mem_dataIn_bits_25(dram1Converter_io_mem_dataIn_bits_25),
    .io_mem_dataIn_bits_26(dram1Converter_io_mem_dataIn_bits_26),
    .io_mem_dataIn_bits_27(dram1Converter_io_mem_dataIn_bits_27),
    .io_mem_dataIn_bits_28(dram1Converter_io_mem_dataIn_bits_28),
    .io_mem_dataIn_bits_29(dram1Converter_io_mem_dataIn_bits_29),
    .io_mem_dataIn_bits_30(dram1Converter_io_mem_dataIn_bits_30),
    .io_mem_dataIn_bits_31(dram1Converter_io_mem_dataIn_bits_31),
    .io_mem_dataOut_ready(dram1Converter_io_mem_dataOut_ready),
    .io_mem_dataOut_valid(dram1Converter_io_mem_dataOut_valid),
    .io_mem_dataOut_bits_0(dram1Converter_io_mem_dataOut_bits_0),
    .io_mem_dataOut_bits_1(dram1Converter_io_mem_dataOut_bits_1),
    .io_mem_dataOut_bits_2(dram1Converter_io_mem_dataOut_bits_2),
    .io_mem_dataOut_bits_3(dram1Converter_io_mem_dataOut_bits_3),
    .io_mem_dataOut_bits_4(dram1Converter_io_mem_dataOut_bits_4),
    .io_mem_dataOut_bits_5(dram1Converter_io_mem_dataOut_bits_5),
    .io_mem_dataOut_bits_6(dram1Converter_io_mem_dataOut_bits_6),
    .io_mem_dataOut_bits_7(dram1Converter_io_mem_dataOut_bits_7),
    .io_mem_dataOut_bits_8(dram1Converter_io_mem_dataOut_bits_8),
    .io_mem_dataOut_bits_9(dram1Converter_io_mem_dataOut_bits_9),
    .io_mem_dataOut_bits_10(dram1Converter_io_mem_dataOut_bits_10),
    .io_mem_dataOut_bits_11(dram1Converter_io_mem_dataOut_bits_11),
    .io_mem_dataOut_bits_12(dram1Converter_io_mem_dataOut_bits_12),
    .io_mem_dataOut_bits_13(dram1Converter_io_mem_dataOut_bits_13),
    .io_mem_dataOut_bits_14(dram1Converter_io_mem_dataOut_bits_14),
    .io_mem_dataOut_bits_15(dram1Converter_io_mem_dataOut_bits_15),
    .io_mem_dataOut_bits_16(dram1Converter_io_mem_dataOut_bits_16),
    .io_mem_dataOut_bits_17(dram1Converter_io_mem_dataOut_bits_17),
    .io_mem_dataOut_bits_18(dram1Converter_io_mem_dataOut_bits_18),
    .io_mem_dataOut_bits_19(dram1Converter_io_mem_dataOut_bits_19),
    .io_mem_dataOut_bits_20(dram1Converter_io_mem_dataOut_bits_20),
    .io_mem_dataOut_bits_21(dram1Converter_io_mem_dataOut_bits_21),
    .io_mem_dataOut_bits_22(dram1Converter_io_mem_dataOut_bits_22),
    .io_mem_dataOut_bits_23(dram1Converter_io_mem_dataOut_bits_23),
    .io_mem_dataOut_bits_24(dram1Converter_io_mem_dataOut_bits_24),
    .io_mem_dataOut_bits_25(dram1Converter_io_mem_dataOut_bits_25),
    .io_mem_dataOut_bits_26(dram1Converter_io_mem_dataOut_bits_26),
    .io_mem_dataOut_bits_27(dram1Converter_io_mem_dataOut_bits_27),
    .io_mem_dataOut_bits_28(dram1Converter_io_mem_dataOut_bits_28),
    .io_mem_dataOut_bits_29(dram1Converter_io_mem_dataOut_bits_29),
    .io_mem_dataOut_bits_30(dram1Converter_io_mem_dataOut_bits_30),
    .io_mem_dataOut_bits_31(dram1Converter_io_mem_dataOut_bits_31),
    .io_axi_writeAddress_ready(dram1Converter_io_axi_writeAddress_ready),
    .io_axi_writeAddress_valid(dram1Converter_io_axi_writeAddress_valid),
    .io_axi_writeAddress_bits_addr(dram1Converter_io_axi_writeAddress_bits_addr),
    .io_axi_writeAddress_bits_len(dram1Converter_io_axi_writeAddress_bits_len),
    .io_axi_writeAddress_bits_cache(dram1Converter_io_axi_writeAddress_bits_cache),
    .io_axi_writeData_ready(dram1Converter_io_axi_writeData_ready),
    .io_axi_writeData_valid(dram1Converter_io_axi_writeData_valid),
    .io_axi_writeData_bits_data(dram1Converter_io_axi_writeData_bits_data),
    .io_axi_writeResponse_ready(dram1Converter_io_axi_writeResponse_ready),
    .io_axi_writeResponse_valid(dram1Converter_io_axi_writeResponse_valid),
    .io_axi_readAddress_ready(dram1Converter_io_axi_readAddress_ready),
    .io_axi_readAddress_valid(dram1Converter_io_axi_readAddress_valid),
    .io_axi_readAddress_bits_addr(dram1Converter_io_axi_readAddress_bits_addr),
    .io_axi_readAddress_bits_len(dram1Converter_io_axi_readAddress_bits_len),
    .io_axi_readAddress_bits_cache(dram1Converter_io_axi_readAddress_bits_cache),
    .io_axi_readData_ready(dram1Converter_io_axi_readData_ready),
    .io_axi_readData_valid(dram1Converter_io_axi_readData_valid),
    .io_axi_readData_bits_data(dram1Converter_io_axi_readData_bits_data),
    .io_axi_readData_bits_last(dram1Converter_io_axi_readData_bits_last),
    .io_addressOffset(dram1Converter_io_addressOffset),
    .io_cacheBehavior(dram1Converter_io_cacheBehavior),
    .io_timeout(dram1Converter_io_timeout),
    .io_tracepoint(dram1Converter_io_tracepoint),
    .io_programCounter(dram1Converter_io_programCounter)
  );
  Queue_45 dram1BoundarySplitter_io_in_q ( // @[Queue.scala 23:19]
    .clock(dram1BoundarySplitter_io_in_q_clock),
    .reset(dram1BoundarySplitter_io_in_q_reset),
    .io_in_writeAddress_ready(dram1BoundarySplitter_io_in_q_io_in_writeAddress_ready),
    .io_in_writeAddress_valid(dram1BoundarySplitter_io_in_q_io_in_writeAddress_valid),
    .io_in_writeAddress_bits_addr(dram1BoundarySplitter_io_in_q_io_in_writeAddress_bits_addr),
    .io_in_writeAddress_bits_len(dram1BoundarySplitter_io_in_q_io_in_writeAddress_bits_len),
    .io_in_writeAddress_bits_cache(dram1BoundarySplitter_io_in_q_io_in_writeAddress_bits_cache),
    .io_in_writeData_ready(dram1BoundarySplitter_io_in_q_io_in_writeData_ready),
    .io_in_writeData_valid(dram1BoundarySplitter_io_in_q_io_in_writeData_valid),
    .io_in_writeData_bits_data(dram1BoundarySplitter_io_in_q_io_in_writeData_bits_data),
    .io_in_writeResponse_ready(dram1BoundarySplitter_io_in_q_io_in_writeResponse_ready),
    .io_in_writeResponse_valid(dram1BoundarySplitter_io_in_q_io_in_writeResponse_valid),
    .io_in_readAddress_ready(dram1BoundarySplitter_io_in_q_io_in_readAddress_ready),
    .io_in_readAddress_valid(dram1BoundarySplitter_io_in_q_io_in_readAddress_valid),
    .io_in_readAddress_bits_addr(dram1BoundarySplitter_io_in_q_io_in_readAddress_bits_addr),
    .io_in_readAddress_bits_len(dram1BoundarySplitter_io_in_q_io_in_readAddress_bits_len),
    .io_in_readAddress_bits_cache(dram1BoundarySplitter_io_in_q_io_in_readAddress_bits_cache),
    .io_in_readData_ready(dram1BoundarySplitter_io_in_q_io_in_readData_ready),
    .io_in_readData_valid(dram1BoundarySplitter_io_in_q_io_in_readData_valid),
    .io_in_readData_bits_data(dram1BoundarySplitter_io_in_q_io_in_readData_bits_data),
    .io_in_readData_bits_last(dram1BoundarySplitter_io_in_q_io_in_readData_bits_last),
    .io_out_writeAddress_ready(dram1BoundarySplitter_io_in_q_io_out_writeAddress_ready),
    .io_out_writeAddress_valid(dram1BoundarySplitter_io_in_q_io_out_writeAddress_valid),
    .io_out_writeAddress_bits_id(dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_id),
    .io_out_writeAddress_bits_addr(dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_addr),
    .io_out_writeAddress_bits_len(dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_len),
    .io_out_writeAddress_bits_size(dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_size),
    .io_out_writeAddress_bits_burst(dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_burst),
    .io_out_writeAddress_bits_lock(dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_lock),
    .io_out_writeAddress_bits_cache(dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_cache),
    .io_out_writeAddress_bits_prot(dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_prot),
    .io_out_writeAddress_bits_qos(dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_qos),
    .io_out_writeData_ready(dram1BoundarySplitter_io_in_q_io_out_writeData_ready),
    .io_out_writeData_valid(dram1BoundarySplitter_io_in_q_io_out_writeData_valid),
    .io_out_writeData_bits_id(dram1BoundarySplitter_io_in_q_io_out_writeData_bits_id),
    .io_out_writeData_bits_data(dram1BoundarySplitter_io_in_q_io_out_writeData_bits_data),
    .io_out_writeData_bits_strb(dram1BoundarySplitter_io_in_q_io_out_writeData_bits_strb),
    .io_out_writeResponse_ready(dram1BoundarySplitter_io_in_q_io_out_writeResponse_ready),
    .io_out_writeResponse_valid(dram1BoundarySplitter_io_in_q_io_out_writeResponse_valid),
    .io_out_readAddress_ready(dram1BoundarySplitter_io_in_q_io_out_readAddress_ready),
    .io_out_readAddress_valid(dram1BoundarySplitter_io_in_q_io_out_readAddress_valid),
    .io_out_readAddress_bits_id(dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_id),
    .io_out_readAddress_bits_addr(dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_addr),
    .io_out_readAddress_bits_len(dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_len),
    .io_out_readAddress_bits_size(dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_size),
    .io_out_readAddress_bits_burst(dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_burst),
    .io_out_readAddress_bits_lock(dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_lock),
    .io_out_readAddress_bits_cache(dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_cache),
    .io_out_readAddress_bits_prot(dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_prot),
    .io_out_readAddress_bits_qos(dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_qos),
    .io_out_readData_ready(dram1BoundarySplitter_io_in_q_io_out_readData_ready),
    .io_out_readData_valid(dram1BoundarySplitter_io_in_q_io_out_readData_valid),
    .io_out_readData_bits_data(dram1BoundarySplitter_io_in_q_io_out_readData_bits_data),
    .io_out_readData_bits_last(dram1BoundarySplitter_io_in_q_io_out_readData_bits_last)
  );
  assign instruction_ready = tcu_io_instruction_ready; // @[AXIWrapperTCU.scala 47:22]
  assign dram0_writeAddress_valid = dram0BoundarySplitter_io_out_writeAddress_valid; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeAddress_bits_id = dram0BoundarySplitter_io_out_writeAddress_bits_id; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeAddress_bits_addr = dram0BoundarySplitter_io_out_writeAddress_bits_addr; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeAddress_bits_len = dram0BoundarySplitter_io_out_writeAddress_bits_len; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeAddress_bits_size = dram0BoundarySplitter_io_out_writeAddress_bits_size; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeAddress_bits_burst = dram0BoundarySplitter_io_out_writeAddress_bits_burst; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeAddress_bits_lock = dram0BoundarySplitter_io_out_writeAddress_bits_lock; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeAddress_bits_cache = dram0BoundarySplitter_io_out_writeAddress_bits_cache; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeAddress_bits_prot = dram0BoundarySplitter_io_out_writeAddress_bits_prot; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeAddress_bits_qos = dram0BoundarySplitter_io_out_writeAddress_bits_qos; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeData_valid = dram0BoundarySplitter_io_out_writeData_valid; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeData_bits_id = dram0BoundarySplitter_io_out_writeData_bits_id; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeData_bits_data = dram0BoundarySplitter_io_out_writeData_bits_data; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeData_bits_strb = dram0BoundarySplitter_io_out_writeData_bits_strb; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeData_bits_last = dram0BoundarySplitter_io_out_writeData_bits_last; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_writeResponse_ready = dram0BoundarySplitter_io_out_writeResponse_ready; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readAddress_valid = dram0BoundarySplitter_io_out_readAddress_valid; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readAddress_bits_id = dram0BoundarySplitter_io_out_readAddress_bits_id; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readAddress_bits_addr = dram0BoundarySplitter_io_out_readAddress_bits_addr; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readAddress_bits_len = dram0BoundarySplitter_io_out_readAddress_bits_len; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readAddress_bits_size = dram0BoundarySplitter_io_out_readAddress_bits_size; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readAddress_bits_burst = dram0BoundarySplitter_io_out_readAddress_bits_burst; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readAddress_bits_lock = dram0BoundarySplitter_io_out_readAddress_bits_lock; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readAddress_bits_cache = dram0BoundarySplitter_io_out_readAddress_bits_cache; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readAddress_bits_prot = dram0BoundarySplitter_io_out_readAddress_bits_prot; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readAddress_bits_qos = dram0BoundarySplitter_io_out_readAddress_bits_qos; // @[AXIWrapperTCU.scala 59:9]
  assign dram0_readData_ready = dram0BoundarySplitter_io_out_readData_ready; // @[AXIWrapperTCU.scala 59:9]
  assign dram1_writeAddress_valid = dram1BoundarySplitter_io_out_writeAddress_valid; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeAddress_bits_id = dram1BoundarySplitter_io_out_writeAddress_bits_id; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeAddress_bits_addr = dram1BoundarySplitter_io_out_writeAddress_bits_addr; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeAddress_bits_len = dram1BoundarySplitter_io_out_writeAddress_bits_len; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeAddress_bits_size = dram1BoundarySplitter_io_out_writeAddress_bits_size; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeAddress_bits_burst = dram1BoundarySplitter_io_out_writeAddress_bits_burst; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeAddress_bits_lock = dram1BoundarySplitter_io_out_writeAddress_bits_lock; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeAddress_bits_cache = dram1BoundarySplitter_io_out_writeAddress_bits_cache; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeAddress_bits_prot = dram1BoundarySplitter_io_out_writeAddress_bits_prot; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeAddress_bits_qos = dram1BoundarySplitter_io_out_writeAddress_bits_qos; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeData_valid = dram1BoundarySplitter_io_out_writeData_valid; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeData_bits_id = dram1BoundarySplitter_io_out_writeData_bits_id; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeData_bits_data = dram1BoundarySplitter_io_out_writeData_bits_data; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeData_bits_strb = dram1BoundarySplitter_io_out_writeData_bits_strb; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeData_bits_last = dram1BoundarySplitter_io_out_writeData_bits_last; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_writeResponse_ready = dram1BoundarySplitter_io_out_writeResponse_ready; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readAddress_valid = dram1BoundarySplitter_io_out_readAddress_valid; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readAddress_bits_id = dram1BoundarySplitter_io_out_readAddress_bits_id; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readAddress_bits_addr = dram1BoundarySplitter_io_out_readAddress_bits_addr; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readAddress_bits_len = dram1BoundarySplitter_io_out_readAddress_bits_len; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readAddress_bits_size = dram1BoundarySplitter_io_out_readAddress_bits_size; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readAddress_bits_burst = dram1BoundarySplitter_io_out_readAddress_bits_burst; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readAddress_bits_lock = dram1BoundarySplitter_io_out_readAddress_bits_lock; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readAddress_bits_cache = dram1BoundarySplitter_io_out_readAddress_bits_cache; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readAddress_bits_prot = dram1BoundarySplitter_io_out_readAddress_bits_prot; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readAddress_bits_qos = dram1BoundarySplitter_io_out_readAddress_bits_qos; // @[AXIWrapperTCU.scala 63:9]
  assign dram1_readData_ready = dram1BoundarySplitter_io_out_readData_ready; // @[AXIWrapperTCU.scala 63:9]
  assign tcu_clock = clock;
  assign tcu_reset = reset;
  assign tcu_io_instruction_valid = instruction_valid; // @[AXIWrapperTCU.scala 47:22]
  assign tcu_io_instruction_bits_opcode = instruction_bits_opcode; // @[AXIWrapperTCU.scala 47:22]
  assign tcu_io_instruction_bits_flags = instruction_bits_flags; // @[AXIWrapperTCU.scala 47:22]
  assign tcu_io_instruction_bits_arguments = instruction_bits_arguments; // @[AXIWrapperTCU.scala 47:22]
  assign tcu_io_dram0_control_ready = dram0Converter_io_mem_control_ready; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_valid = dram0Converter_io_mem_dataIn_valid; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_0 = dram0Converter_io_mem_dataIn_bits_0; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_1 = dram0Converter_io_mem_dataIn_bits_1; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_2 = dram0Converter_io_mem_dataIn_bits_2; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_3 = dram0Converter_io_mem_dataIn_bits_3; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_4 = dram0Converter_io_mem_dataIn_bits_4; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_5 = dram0Converter_io_mem_dataIn_bits_5; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_6 = dram0Converter_io_mem_dataIn_bits_6; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_7 = dram0Converter_io_mem_dataIn_bits_7; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_8 = dram0Converter_io_mem_dataIn_bits_8; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_9 = dram0Converter_io_mem_dataIn_bits_9; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_10 = dram0Converter_io_mem_dataIn_bits_10; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_11 = dram0Converter_io_mem_dataIn_bits_11; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_12 = dram0Converter_io_mem_dataIn_bits_12; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_13 = dram0Converter_io_mem_dataIn_bits_13; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_14 = dram0Converter_io_mem_dataIn_bits_14; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_15 = dram0Converter_io_mem_dataIn_bits_15; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_16 = dram0Converter_io_mem_dataIn_bits_16; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_17 = dram0Converter_io_mem_dataIn_bits_17; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_18 = dram0Converter_io_mem_dataIn_bits_18; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_19 = dram0Converter_io_mem_dataIn_bits_19; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_20 = dram0Converter_io_mem_dataIn_bits_20; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_21 = dram0Converter_io_mem_dataIn_bits_21; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_22 = dram0Converter_io_mem_dataIn_bits_22; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_23 = dram0Converter_io_mem_dataIn_bits_23; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_24 = dram0Converter_io_mem_dataIn_bits_24; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_25 = dram0Converter_io_mem_dataIn_bits_25; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_26 = dram0Converter_io_mem_dataIn_bits_26; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_27 = dram0Converter_io_mem_dataIn_bits_27; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_28 = dram0Converter_io_mem_dataIn_bits_28; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_29 = dram0Converter_io_mem_dataIn_bits_29; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_30 = dram0Converter_io_mem_dataIn_bits_30; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataIn_bits_31 = dram0Converter_io_mem_dataIn_bits_31; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram0_dataOut_ready = dram0Converter_io_mem_dataOut_ready; // @[AXIWrapperTCU.scala 75:25]
  assign tcu_io_dram1_control_ready = dram1Converter_io_mem_control_ready; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_valid = dram1Converter_io_mem_dataIn_valid; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_0 = dram1Converter_io_mem_dataIn_bits_0; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_1 = dram1Converter_io_mem_dataIn_bits_1; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_2 = dram1Converter_io_mem_dataIn_bits_2; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_3 = dram1Converter_io_mem_dataIn_bits_3; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_4 = dram1Converter_io_mem_dataIn_bits_4; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_5 = dram1Converter_io_mem_dataIn_bits_5; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_6 = dram1Converter_io_mem_dataIn_bits_6; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_7 = dram1Converter_io_mem_dataIn_bits_7; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_8 = dram1Converter_io_mem_dataIn_bits_8; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_9 = dram1Converter_io_mem_dataIn_bits_9; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_10 = dram1Converter_io_mem_dataIn_bits_10; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_11 = dram1Converter_io_mem_dataIn_bits_11; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_12 = dram1Converter_io_mem_dataIn_bits_12; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_13 = dram1Converter_io_mem_dataIn_bits_13; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_14 = dram1Converter_io_mem_dataIn_bits_14; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_15 = dram1Converter_io_mem_dataIn_bits_15; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_16 = dram1Converter_io_mem_dataIn_bits_16; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_17 = dram1Converter_io_mem_dataIn_bits_17; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_18 = dram1Converter_io_mem_dataIn_bits_18; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_19 = dram1Converter_io_mem_dataIn_bits_19; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_20 = dram1Converter_io_mem_dataIn_bits_20; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_21 = dram1Converter_io_mem_dataIn_bits_21; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_22 = dram1Converter_io_mem_dataIn_bits_22; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_23 = dram1Converter_io_mem_dataIn_bits_23; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_24 = dram1Converter_io_mem_dataIn_bits_24; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_25 = dram1Converter_io_mem_dataIn_bits_25; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_26 = dram1Converter_io_mem_dataIn_bits_26; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_27 = dram1Converter_io_mem_dataIn_bits_27; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_28 = dram1Converter_io_mem_dataIn_bits_28; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_29 = dram1Converter_io_mem_dataIn_bits_29; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_30 = dram1Converter_io_mem_dataIn_bits_30; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataIn_bits_31 = dram1Converter_io_mem_dataIn_bits_31; // @[AXIWrapperTCU.scala 92:25]
  assign tcu_io_dram1_dataOut_ready = dram1Converter_io_mem_dataOut_ready; // @[AXIWrapperTCU.scala 92:25]
  assign dram0BoundarySplitter_clock = clock;
  assign dram0BoundarySplitter_reset = reset;
  assign dram0BoundarySplitter_io_in_writeAddress_valid = dram0BoundarySplitter_io_in_q_io_out_writeAddress_valid; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeAddress_bits_id = dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_id; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeAddress_bits_addr =
    dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_addr; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeAddress_bits_len = dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_len; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeAddress_bits_size =
    dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_size; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeAddress_bits_burst =
    dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_burst; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeAddress_bits_lock =
    dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_lock; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeAddress_bits_cache =
    dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_cache; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeAddress_bits_prot =
    dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_prot; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeAddress_bits_qos = dram0BoundarySplitter_io_in_q_io_out_writeAddress_bits_qos; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeData_valid = dram0BoundarySplitter_io_in_q_io_out_writeData_valid; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeData_bits_id = dram0BoundarySplitter_io_in_q_io_out_writeData_bits_id; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeData_bits_data = dram0BoundarySplitter_io_in_q_io_out_writeData_bits_data; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeData_bits_strb = dram0BoundarySplitter_io_in_q_io_out_writeData_bits_strb; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_writeResponse_ready = dram0BoundarySplitter_io_in_q_io_out_writeResponse_ready; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readAddress_valid = dram0BoundarySplitter_io_in_q_io_out_readAddress_valid; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readAddress_bits_id = dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_id; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readAddress_bits_addr = dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_addr; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readAddress_bits_len = dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_len; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readAddress_bits_size = dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_size; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readAddress_bits_burst =
    dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_burst; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readAddress_bits_lock = dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_lock; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readAddress_bits_cache =
    dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_cache; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readAddress_bits_prot = dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_prot; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readAddress_bits_qos = dram0BoundarySplitter_io_in_q_io_out_readAddress_bits_qos; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_readData_ready = dram0BoundarySplitter_io_in_q_io_out_readData_ready; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_out_writeAddress_ready = dram0_writeAddress_ready; // @[AXIWrapperTCU.scala 59:9]
  assign dram0BoundarySplitter_io_out_writeData_ready = dram0_writeData_ready; // @[AXIWrapperTCU.scala 59:9]
  assign dram0BoundarySplitter_io_out_writeResponse_valid = dram0_writeResponse_valid; // @[AXIWrapperTCU.scala 59:9]
  assign dram0BoundarySplitter_io_out_readAddress_ready = dram0_readAddress_ready; // @[AXIWrapperTCU.scala 59:9]
  assign dram0BoundarySplitter_io_out_readData_valid = dram0_readData_valid; // @[AXIWrapperTCU.scala 59:9]
  assign dram0BoundarySplitter_io_out_readData_bits_data = dram0_readData_bits_data; // @[AXIWrapperTCU.scala 59:9]
  assign dram1BoundarySplitter_clock = clock;
  assign dram1BoundarySplitter_reset = reset;
  assign dram1BoundarySplitter_io_in_writeAddress_valid = dram1BoundarySplitter_io_in_q_io_out_writeAddress_valid; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeAddress_bits_id = dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_id; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeAddress_bits_addr =
    dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_addr; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeAddress_bits_len = dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_len; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeAddress_bits_size =
    dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_size; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeAddress_bits_burst =
    dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_burst; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeAddress_bits_lock =
    dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_lock; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeAddress_bits_cache =
    dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_cache; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeAddress_bits_prot =
    dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_prot; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeAddress_bits_qos = dram1BoundarySplitter_io_in_q_io_out_writeAddress_bits_qos; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeData_valid = dram1BoundarySplitter_io_in_q_io_out_writeData_valid; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeData_bits_id = dram1BoundarySplitter_io_in_q_io_out_writeData_bits_id; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeData_bits_data = dram1BoundarySplitter_io_in_q_io_out_writeData_bits_data; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeData_bits_strb = dram1BoundarySplitter_io_in_q_io_out_writeData_bits_strb; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_writeResponse_ready = dram1BoundarySplitter_io_in_q_io_out_writeResponse_ready; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readAddress_valid = dram1BoundarySplitter_io_in_q_io_out_readAddress_valid; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readAddress_bits_id = dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_id; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readAddress_bits_addr = dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_addr; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readAddress_bits_len = dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_len; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readAddress_bits_size = dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_size; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readAddress_bits_burst =
    dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_burst; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readAddress_bits_lock = dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_lock; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readAddress_bits_cache =
    dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_cache; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readAddress_bits_prot = dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_prot; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readAddress_bits_qos = dram1BoundarySplitter_io_in_q_io_out_readAddress_bits_qos; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_readData_ready = dram1BoundarySplitter_io_in_q_io_out_readData_ready; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_out_writeAddress_ready = dram1_writeAddress_ready; // @[AXIWrapperTCU.scala 63:9]
  assign dram1BoundarySplitter_io_out_writeData_ready = dram1_writeData_ready; // @[AXIWrapperTCU.scala 63:9]
  assign dram1BoundarySplitter_io_out_writeResponse_valid = dram1_writeResponse_valid; // @[AXIWrapperTCU.scala 63:9]
  assign dram1BoundarySplitter_io_out_readAddress_ready = dram1_readAddress_ready; // @[AXIWrapperTCU.scala 63:9]
  assign dram1BoundarySplitter_io_out_readData_valid = dram1_readData_valid; // @[AXIWrapperTCU.scala 63:9]
  assign dram1BoundarySplitter_io_out_readData_bits_data = dram1_readData_bits_data; // @[AXIWrapperTCU.scala 63:9]
  assign dram0Converter_clock = clock;
  assign dram0Converter_reset = reset;
  assign dram0Converter_io_mem_control_valid = tcu_io_dram0_control_valid; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_control_bits_write = tcu_io_dram0_control_bits_write; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_control_bits_address = tcu_io_dram0_control_bits_address; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_control_bits_size = tcu_io_dram0_control_bits_size; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataIn_ready = tcu_io_dram0_dataIn_ready; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_valid = tcu_io_dram0_dataOut_valid; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_0 = tcu_io_dram0_dataOut_bits_0; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_1 = tcu_io_dram0_dataOut_bits_1; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_2 = tcu_io_dram0_dataOut_bits_2; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_3 = tcu_io_dram0_dataOut_bits_3; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_4 = tcu_io_dram0_dataOut_bits_4; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_5 = tcu_io_dram0_dataOut_bits_5; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_6 = tcu_io_dram0_dataOut_bits_6; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_7 = tcu_io_dram0_dataOut_bits_7; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_8 = tcu_io_dram0_dataOut_bits_8; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_9 = tcu_io_dram0_dataOut_bits_9; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_10 = tcu_io_dram0_dataOut_bits_10; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_11 = tcu_io_dram0_dataOut_bits_11; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_12 = tcu_io_dram0_dataOut_bits_12; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_13 = tcu_io_dram0_dataOut_bits_13; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_14 = tcu_io_dram0_dataOut_bits_14; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_15 = tcu_io_dram0_dataOut_bits_15; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_16 = tcu_io_dram0_dataOut_bits_16; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_17 = tcu_io_dram0_dataOut_bits_17; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_18 = tcu_io_dram0_dataOut_bits_18; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_19 = tcu_io_dram0_dataOut_bits_19; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_20 = tcu_io_dram0_dataOut_bits_20; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_21 = tcu_io_dram0_dataOut_bits_21; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_22 = tcu_io_dram0_dataOut_bits_22; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_23 = tcu_io_dram0_dataOut_bits_23; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_24 = tcu_io_dram0_dataOut_bits_24; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_25 = tcu_io_dram0_dataOut_bits_25; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_26 = tcu_io_dram0_dataOut_bits_26; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_27 = tcu_io_dram0_dataOut_bits_27; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_28 = tcu_io_dram0_dataOut_bits_28; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_29 = tcu_io_dram0_dataOut_bits_29; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_30 = tcu_io_dram0_dataOut_bits_30; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_mem_dataOut_bits_31 = tcu_io_dram0_dataOut_bits_31; // @[AXIWrapperTCU.scala 75:25]
  assign dram0Converter_io_axi_writeAddress_ready = dram0BoundarySplitter_io_in_q_io_in_writeAddress_ready; // @[Queue.scala 24:13]
  assign dram0Converter_io_axi_writeData_ready = dram0BoundarySplitter_io_in_q_io_in_writeData_ready; // @[Queue.scala 24:13]
  assign dram0Converter_io_axi_writeResponse_valid = dram0BoundarySplitter_io_in_q_io_in_writeResponse_valid; // @[Queue.scala 24:13]
  assign dram0Converter_io_axi_readAddress_ready = dram0BoundarySplitter_io_in_q_io_in_readAddress_ready; // @[Queue.scala 24:13]
  assign dram0Converter_io_axi_readData_valid = dram0BoundarySplitter_io_in_q_io_in_readData_valid; // @[Queue.scala 24:13]
  assign dram0Converter_io_axi_readData_bits_data = dram0BoundarySplitter_io_in_q_io_in_readData_bits_data; // @[Queue.scala 24:13]
  assign dram0Converter_io_axi_readData_bits_last = dram0BoundarySplitter_io_in_q_io_in_readData_bits_last; // @[Queue.scala 24:13]
  assign dram0Converter_io_addressOffset = tcu_io_config_dram0AddressOffset; // @[AXIWrapperTCU.scala 76:35]
  assign dram0Converter_io_cacheBehavior = tcu_io_config_dram0CacheBehaviour; // @[AXIWrapperTCU.scala 77:35]
  assign dram0Converter_io_timeout = tcu_io_timeout; // @[AXIWrapperTCU.scala 78:29]
  assign dram0Converter_io_tracepoint = tcu_io_tracepoint; // @[AXIWrapperTCU.scala 79:32]
  assign dram0Converter_io_programCounter = tcu_io_programCounter; // @[AXIWrapperTCU.scala 80:36]
  assign dram0BoundarySplitter_io_in_q_clock = clock;
  assign dram0BoundarySplitter_io_in_q_reset = reset;
  assign dram0BoundarySplitter_io_in_q_io_in_writeAddress_valid = dram0Converter_io_axi_writeAddress_valid; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_writeAddress_bits_addr = dram0Converter_io_axi_writeAddress_bits_addr; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_writeAddress_bits_len = dram0Converter_io_axi_writeAddress_bits_len; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_writeAddress_bits_cache = dram0Converter_io_axi_writeAddress_bits_cache; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_writeData_valid = dram0Converter_io_axi_writeData_valid; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_writeData_bits_data = dram0Converter_io_axi_writeData_bits_data; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_writeResponse_ready = dram0Converter_io_axi_writeResponse_ready; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_readAddress_valid = dram0Converter_io_axi_readAddress_valid; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_readAddress_bits_addr = dram0Converter_io_axi_readAddress_bits_addr; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_readAddress_bits_len = dram0Converter_io_axi_readAddress_bits_len; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_readAddress_bits_cache = dram0Converter_io_axi_readAddress_bits_cache; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_in_readData_ready = dram0Converter_io_axi_readData_ready; // @[Queue.scala 24:13]
  assign dram0BoundarySplitter_io_in_q_io_out_writeAddress_ready = dram0BoundarySplitter_io_in_writeAddress_ready; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_q_io_out_writeData_ready = dram0BoundarySplitter_io_in_writeData_ready; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_q_io_out_writeResponse_valid = dram0BoundarySplitter_io_in_writeResponse_valid; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_q_io_out_readAddress_ready = dram0BoundarySplitter_io_in_readAddress_ready; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_q_io_out_readData_valid = dram0BoundarySplitter_io_in_readData_valid; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_q_io_out_readData_bits_data = dram0BoundarySplitter_io_in_readData_bits_data; // @[AXIWrapperTCU.scala 74:31]
  assign dram0BoundarySplitter_io_in_q_io_out_readData_bits_last = dram0BoundarySplitter_io_in_readData_bits_last; // @[AXIWrapperTCU.scala 74:31]
  assign dram1Converter_clock = clock;
  assign dram1Converter_reset = reset;
  assign dram1Converter_io_mem_control_valid = tcu_io_dram1_control_valid; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_control_bits_write = tcu_io_dram1_control_bits_write; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_control_bits_address = tcu_io_dram1_control_bits_address; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_control_bits_size = tcu_io_dram1_control_bits_size; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataIn_ready = tcu_io_dram1_dataIn_ready; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_valid = tcu_io_dram1_dataOut_valid; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_0 = tcu_io_dram1_dataOut_bits_0; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_1 = tcu_io_dram1_dataOut_bits_1; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_2 = tcu_io_dram1_dataOut_bits_2; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_3 = tcu_io_dram1_dataOut_bits_3; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_4 = tcu_io_dram1_dataOut_bits_4; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_5 = tcu_io_dram1_dataOut_bits_5; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_6 = tcu_io_dram1_dataOut_bits_6; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_7 = tcu_io_dram1_dataOut_bits_7; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_8 = tcu_io_dram1_dataOut_bits_8; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_9 = tcu_io_dram1_dataOut_bits_9; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_10 = tcu_io_dram1_dataOut_bits_10; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_11 = tcu_io_dram1_dataOut_bits_11; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_12 = tcu_io_dram1_dataOut_bits_12; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_13 = tcu_io_dram1_dataOut_bits_13; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_14 = tcu_io_dram1_dataOut_bits_14; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_15 = tcu_io_dram1_dataOut_bits_15; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_16 = tcu_io_dram1_dataOut_bits_16; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_17 = tcu_io_dram1_dataOut_bits_17; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_18 = tcu_io_dram1_dataOut_bits_18; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_19 = tcu_io_dram1_dataOut_bits_19; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_20 = tcu_io_dram1_dataOut_bits_20; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_21 = tcu_io_dram1_dataOut_bits_21; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_22 = tcu_io_dram1_dataOut_bits_22; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_23 = tcu_io_dram1_dataOut_bits_23; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_24 = tcu_io_dram1_dataOut_bits_24; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_25 = tcu_io_dram1_dataOut_bits_25; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_26 = tcu_io_dram1_dataOut_bits_26; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_27 = tcu_io_dram1_dataOut_bits_27; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_28 = tcu_io_dram1_dataOut_bits_28; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_29 = tcu_io_dram1_dataOut_bits_29; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_30 = tcu_io_dram1_dataOut_bits_30; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_mem_dataOut_bits_31 = tcu_io_dram1_dataOut_bits_31; // @[AXIWrapperTCU.scala 92:25]
  assign dram1Converter_io_axi_writeAddress_ready = dram1BoundarySplitter_io_in_q_io_in_writeAddress_ready; // @[Queue.scala 24:13]
  assign dram1Converter_io_axi_writeData_ready = dram1BoundarySplitter_io_in_q_io_in_writeData_ready; // @[Queue.scala 24:13]
  assign dram1Converter_io_axi_writeResponse_valid = dram1BoundarySplitter_io_in_q_io_in_writeResponse_valid; // @[Queue.scala 24:13]
  assign dram1Converter_io_axi_readAddress_ready = dram1BoundarySplitter_io_in_q_io_in_readAddress_ready; // @[Queue.scala 24:13]
  assign dram1Converter_io_axi_readData_valid = dram1BoundarySplitter_io_in_q_io_in_readData_valid; // @[Queue.scala 24:13]
  assign dram1Converter_io_axi_readData_bits_data = dram1BoundarySplitter_io_in_q_io_in_readData_bits_data; // @[Queue.scala 24:13]
  assign dram1Converter_io_axi_readData_bits_last = dram1BoundarySplitter_io_in_q_io_in_readData_bits_last; // @[Queue.scala 24:13]
  assign dram1Converter_io_addressOffset = tcu_io_config_dram1AddressOffset; // @[AXIWrapperTCU.scala 93:35]
  assign dram1Converter_io_cacheBehavior = tcu_io_config_dram1CacheBehaviour; // @[AXIWrapperTCU.scala 94:35]
  assign dram1Converter_io_timeout = tcu_io_timeout; // @[AXIWrapperTCU.scala 95:29]
  assign dram1Converter_io_tracepoint = tcu_io_tracepoint; // @[AXIWrapperTCU.scala 96:32]
  assign dram1Converter_io_programCounter = tcu_io_programCounter; // @[AXIWrapperTCU.scala 97:36]
  assign dram1BoundarySplitter_io_in_q_clock = clock;
  assign dram1BoundarySplitter_io_in_q_reset = reset;
  assign dram1BoundarySplitter_io_in_q_io_in_writeAddress_valid = dram1Converter_io_axi_writeAddress_valid; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_writeAddress_bits_addr = dram1Converter_io_axi_writeAddress_bits_addr; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_writeAddress_bits_len = dram1Converter_io_axi_writeAddress_bits_len; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_writeAddress_bits_cache = dram1Converter_io_axi_writeAddress_bits_cache; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_writeData_valid = dram1Converter_io_axi_writeData_valid; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_writeData_bits_data = dram1Converter_io_axi_writeData_bits_data; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_writeResponse_ready = dram1Converter_io_axi_writeResponse_ready; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_readAddress_valid = dram1Converter_io_axi_readAddress_valid; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_readAddress_bits_addr = dram1Converter_io_axi_readAddress_bits_addr; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_readAddress_bits_len = dram1Converter_io_axi_readAddress_bits_len; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_readAddress_bits_cache = dram1Converter_io_axi_readAddress_bits_cache; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_in_readData_ready = dram1Converter_io_axi_readData_ready; // @[Queue.scala 24:13]
  assign dram1BoundarySplitter_io_in_q_io_out_writeAddress_ready = dram1BoundarySplitter_io_in_writeAddress_ready; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_q_io_out_writeData_ready = dram1BoundarySplitter_io_in_writeData_ready; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_q_io_out_writeResponse_valid = dram1BoundarySplitter_io_in_writeResponse_valid; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_q_io_out_readAddress_ready = dram1BoundarySplitter_io_in_readAddress_ready; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_q_io_out_readData_valid = dram1BoundarySplitter_io_in_readData_valid; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_q_io_out_readData_bits_data = dram1BoundarySplitter_io_in_readData_bits_data; // @[AXIWrapperTCU.scala 91:31]
  assign dram1BoundarySplitter_io_in_q_io_out_readData_bits_last = dram1BoundarySplitter_io_in_readData_bits_last; // @[AXIWrapperTCU.scala 91:31]
endmodule
module WidthConverter(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits,
  input          io_out_ready,
  output         io_out_valid,
  output [71:0]  io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] arr_0; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_1; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_2; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_3; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_4; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_5; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_6; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_7; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_8; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_9; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_10; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_11; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_12; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_13; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_14; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_15; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_16; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_17; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_18; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_19; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_20; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_21; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_22; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_23; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_24; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_25; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_26; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_27; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_28; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_29; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_30; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_31; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_32; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_33; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_34; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_35; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_36; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_37; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_38; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_39; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_40; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_41; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_42; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_43; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_44; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_45; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_46; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_47; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_48; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_49; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_50; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_51; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_52; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_53; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_54; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_55; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_56; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_57; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_58; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_59; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_60; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_61; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_62; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_63; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_64; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_65; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_66; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_67; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_68; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_69; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_70; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_71; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_72; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_73; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_74; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_75; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_76; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_77; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_78; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_79; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_80; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_81; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_82; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_83; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_84; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_85; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_86; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_87; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_88; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_89; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_90; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_91; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_92; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_93; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_94; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_95; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_96; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_97; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_98; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_99; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_100; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_101; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_102; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_103; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_104; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_105; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_106; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_107; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_108; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_109; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_110; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_111; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_112; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_113; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_114; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_115; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_116; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_117; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_118; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_119; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_120; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_121; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_122; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_123; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_124; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_125; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_126; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_127; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_128; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_129; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_130; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_131; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_132; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_133; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_134; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_135; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_136; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_137; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_138; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_139; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_140; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_141; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_142; // @[WidthConverter.scala 24:29]
  reg [7:0] arr_143; // @[WidthConverter.scala 24:29]
  reg [7:0] enqPtr; // @[WidthConverter.scala 25:29]
  reg [7:0] deqPtr; // @[WidthConverter.scala 26:29]
  reg  maybeFull; // @[WidthConverter.scala 27:29]
  wire  doEnq = io_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
  wire  doDeq = io_out_ready & io_out_valid; // @[Decoupled.scala 50:35]
  wire  ptrMatch = enqPtr == deqPtr; // @[WidthConverter.scala 30:29]
  wire [8:0] enqPtrNext = enqPtr + 8'h10; // @[WidthConverter.scala 31:29]
  wire [8:0] deqPtrNext = deqPtr + 8'h9; // @[WidthConverter.scala 32:29]
  wire  _full_T = enqPtr < deqPtr; // @[WidthConverter.scala 38:18]
  wire [8:0] _GEN_3747 = {{1'd0}, deqPtr}; // @[WidthConverter.scala 39:22]
  wire  _full_T_1 = enqPtrNext > _GEN_3747; // @[WidthConverter.scala 39:22]
  wire  _full_T_2 = enqPtrNext > 9'h90; // @[WidthConverter.scala 41:24]
  wire [8:0] _GEN_3749 = enqPtrNext % 9'h90; // @[WidthConverter.scala 42:25]
  wire  _full_T_4 = _GEN_3749[7:0] > deqPtr; // @[WidthConverter.scala 42:40]
  wire  _full_T_5 = _full_T_2 & _full_T_4; // @[WidthConverter.scala 40:22]
  wire  _full_T_6 = _full_T ? _full_T_1 : _full_T_5; // @[WidthConverter.scala 37:20]
  wire  full = ptrMatch ? maybeFull : _full_T_6; // @[WidthConverter.scala 34:18]
  wire  _empty_T = ~maybeFull; // @[WidthConverter.scala 49:7]
  wire  _empty_T_1 = deqPtr < enqPtr; // @[WidthConverter.scala 51:16]
  wire [8:0] _GEN_3748 = {{1'd0}, enqPtr}; // @[WidthConverter.scala 52:20]
  wire  _empty_T_2 = deqPtrNext > _GEN_3748; // @[WidthConverter.scala 52:20]
  wire  _empty_T_3 = deqPtrNext > 9'h90; // @[WidthConverter.scala 54:22]
  wire [8:0] _GEN_3750 = deqPtrNext % 9'h90; // @[WidthConverter.scala 55:23]
  wire  _empty_T_5 = _GEN_3750[7:0] > enqPtr; // @[WidthConverter.scala 55:38]
  wire  _empty_T_6 = _empty_T_3 & _empty_T_5; // @[WidthConverter.scala 53:20]
  wire  _empty_T_7 = _empty_T_1 ? _empty_T_2 : _empty_T_6; // @[WidthConverter.scala 50:18]
  wire  empty = ptrMatch ? _empty_T : _empty_T_7; // @[WidthConverter.scala 47:28]
  wire [7:0] _GEN_1 = 8'h0 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_0; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_2 = 8'h1 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_1; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_3 = 8'h2 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_2; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_4 = 8'h3 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_3; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_5 = 8'h4 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_4; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_6 = 8'h5 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_5; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_7 = 8'h6 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_6; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_8 = 8'h7 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_7; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_9 = 8'h8 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_8; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_10 = 8'h9 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_9; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_11 = 8'ha == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_10; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_12 = 8'hb == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_11; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_13 = 8'hc == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_12; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_14 = 8'hd == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_13; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_15 = 8'he == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_14; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_16 = 8'hf == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_15; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_17 = 8'h10 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_16; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_18 = 8'h11 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_17; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_19 = 8'h12 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_18; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_20 = 8'h13 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_19; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_21 = 8'h14 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_20; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_22 = 8'h15 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_21; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_23 = 8'h16 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_22; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_24 = 8'h17 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_23; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_25 = 8'h18 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_24; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_26 = 8'h19 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_25; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_27 = 8'h1a == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_26; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_28 = 8'h1b == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_27; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_29 = 8'h1c == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_28; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_30 = 8'h1d == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_29; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_31 = 8'h1e == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_30; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_32 = 8'h1f == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_31; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_33 = 8'h20 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_32; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_34 = 8'h21 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_33; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_35 = 8'h22 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_34; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_36 = 8'h23 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_35; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_37 = 8'h24 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_36; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_38 = 8'h25 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_37; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_39 = 8'h26 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_38; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_40 = 8'h27 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_39; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_41 = 8'h28 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_40; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_42 = 8'h29 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_41; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_43 = 8'h2a == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_42; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_44 = 8'h2b == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_43; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_45 = 8'h2c == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_44; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_46 = 8'h2d == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_45; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_47 = 8'h2e == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_46; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_48 = 8'h2f == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_47; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_49 = 8'h30 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_48; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_50 = 8'h31 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_49; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_51 = 8'h32 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_50; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_52 = 8'h33 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_51; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_53 = 8'h34 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_52; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_54 = 8'h35 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_53; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_55 = 8'h36 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_54; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_56 = 8'h37 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_55; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_57 = 8'h38 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_56; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_58 = 8'h39 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_57; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_59 = 8'h3a == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_58; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_60 = 8'h3b == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_59; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_61 = 8'h3c == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_60; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_62 = 8'h3d == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_61; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_63 = 8'h3e == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_62; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_64 = 8'h3f == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_63; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_65 = 8'h40 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_64; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_66 = 8'h41 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_65; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_67 = 8'h42 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_66; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_68 = 8'h43 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_67; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_69 = 8'h44 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_68; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_70 = 8'h45 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_69; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_71 = 8'h46 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_70; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_72 = 8'h47 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_71; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_73 = 8'h48 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_72; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_74 = 8'h49 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_73; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_75 = 8'h4a == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_74; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_76 = 8'h4b == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_75; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_77 = 8'h4c == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_76; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_78 = 8'h4d == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_77; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_79 = 8'h4e == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_78; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_80 = 8'h4f == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_79; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_81 = 8'h50 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_80; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_82 = 8'h51 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_81; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_83 = 8'h52 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_82; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_84 = 8'h53 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_83; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_85 = 8'h54 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_84; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_86 = 8'h55 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_85; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_87 = 8'h56 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_86; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_88 = 8'h57 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_87; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_89 = 8'h58 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_88; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_90 = 8'h59 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_89; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_91 = 8'h5a == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_90; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_92 = 8'h5b == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_91; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_93 = 8'h5c == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_92; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_94 = 8'h5d == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_93; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_95 = 8'h5e == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_94; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_96 = 8'h5f == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_95; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_97 = 8'h60 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_96; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_98 = 8'h61 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_97; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_99 = 8'h62 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_98; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_100 = 8'h63 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_99; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_101 = 8'h64 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_100; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_102 = 8'h65 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_101; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_103 = 8'h66 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_102; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_104 = 8'h67 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_103; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_105 = 8'h68 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_104; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_106 = 8'h69 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_105; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_107 = 8'h6a == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_106; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_108 = 8'h6b == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_107; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_109 = 8'h6c == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_108; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_110 = 8'h6d == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_109; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_111 = 8'h6e == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_110; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_112 = 8'h6f == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_111; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_113 = 8'h70 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_112; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_114 = 8'h71 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_113; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_115 = 8'h72 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_114; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_116 = 8'h73 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_115; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_117 = 8'h74 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_116; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_118 = 8'h75 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_117; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_119 = 8'h76 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_118; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_120 = 8'h77 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_119; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_121 = 8'h78 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_120; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_122 = 8'h79 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_121; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_123 = 8'h7a == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_122; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_124 = 8'h7b == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_123; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_125 = 8'h7c == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_124; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_126 = 8'h7d == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_125; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_127 = 8'h7e == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_126; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_128 = 8'h7f == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_127; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_129 = 8'h80 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_128; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_130 = 8'h81 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_129; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_131 = 8'h82 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_130; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_132 = 8'h83 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_131; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_133 = 8'h84 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_132; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_134 = 8'h85 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_133; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_135 = 8'h86 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_134; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_136 = 8'h87 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_135; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_137 = 8'h88 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_136; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_138 = 8'h89 == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_137; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_139 = 8'h8a == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_138; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_140 = 8'h8b == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_139; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_141 = 8'h8c == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_140; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_142 = 8'h8d == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_141; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_143 = 8'h8e == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_142; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _GEN_144 = 8'h8f == _GEN_3748[7:0] ? io_in_bits[7:0] : arr_143; // @[WidthConverter.scala 67:{27,27} 24:29]
  wire [7:0] _T_4 = enqPtr + 8'h1; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_145 = 8'h0 == _T_4 ? io_in_bits[15:8] : _GEN_1; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_146 = 8'h1 == _T_4 ? io_in_bits[15:8] : _GEN_2; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_147 = 8'h2 == _T_4 ? io_in_bits[15:8] : _GEN_3; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_148 = 8'h3 == _T_4 ? io_in_bits[15:8] : _GEN_4; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_149 = 8'h4 == _T_4 ? io_in_bits[15:8] : _GEN_5; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_150 = 8'h5 == _T_4 ? io_in_bits[15:8] : _GEN_6; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_151 = 8'h6 == _T_4 ? io_in_bits[15:8] : _GEN_7; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_152 = 8'h7 == _T_4 ? io_in_bits[15:8] : _GEN_8; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_153 = 8'h8 == _T_4 ? io_in_bits[15:8] : _GEN_9; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_154 = 8'h9 == _T_4 ? io_in_bits[15:8] : _GEN_10; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_155 = 8'ha == _T_4 ? io_in_bits[15:8] : _GEN_11; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_156 = 8'hb == _T_4 ? io_in_bits[15:8] : _GEN_12; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_157 = 8'hc == _T_4 ? io_in_bits[15:8] : _GEN_13; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_158 = 8'hd == _T_4 ? io_in_bits[15:8] : _GEN_14; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_159 = 8'he == _T_4 ? io_in_bits[15:8] : _GEN_15; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_160 = 8'hf == _T_4 ? io_in_bits[15:8] : _GEN_16; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_161 = 8'h10 == _T_4 ? io_in_bits[15:8] : _GEN_17; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_162 = 8'h11 == _T_4 ? io_in_bits[15:8] : _GEN_18; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_163 = 8'h12 == _T_4 ? io_in_bits[15:8] : _GEN_19; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_164 = 8'h13 == _T_4 ? io_in_bits[15:8] : _GEN_20; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_165 = 8'h14 == _T_4 ? io_in_bits[15:8] : _GEN_21; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_166 = 8'h15 == _T_4 ? io_in_bits[15:8] : _GEN_22; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_167 = 8'h16 == _T_4 ? io_in_bits[15:8] : _GEN_23; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_168 = 8'h17 == _T_4 ? io_in_bits[15:8] : _GEN_24; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_169 = 8'h18 == _T_4 ? io_in_bits[15:8] : _GEN_25; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_170 = 8'h19 == _T_4 ? io_in_bits[15:8] : _GEN_26; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_171 = 8'h1a == _T_4 ? io_in_bits[15:8] : _GEN_27; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_172 = 8'h1b == _T_4 ? io_in_bits[15:8] : _GEN_28; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_173 = 8'h1c == _T_4 ? io_in_bits[15:8] : _GEN_29; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_174 = 8'h1d == _T_4 ? io_in_bits[15:8] : _GEN_30; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_175 = 8'h1e == _T_4 ? io_in_bits[15:8] : _GEN_31; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_176 = 8'h1f == _T_4 ? io_in_bits[15:8] : _GEN_32; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_177 = 8'h20 == _T_4 ? io_in_bits[15:8] : _GEN_33; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_178 = 8'h21 == _T_4 ? io_in_bits[15:8] : _GEN_34; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_179 = 8'h22 == _T_4 ? io_in_bits[15:8] : _GEN_35; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_180 = 8'h23 == _T_4 ? io_in_bits[15:8] : _GEN_36; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_181 = 8'h24 == _T_4 ? io_in_bits[15:8] : _GEN_37; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_182 = 8'h25 == _T_4 ? io_in_bits[15:8] : _GEN_38; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_183 = 8'h26 == _T_4 ? io_in_bits[15:8] : _GEN_39; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_184 = 8'h27 == _T_4 ? io_in_bits[15:8] : _GEN_40; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_185 = 8'h28 == _T_4 ? io_in_bits[15:8] : _GEN_41; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_186 = 8'h29 == _T_4 ? io_in_bits[15:8] : _GEN_42; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_187 = 8'h2a == _T_4 ? io_in_bits[15:8] : _GEN_43; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_188 = 8'h2b == _T_4 ? io_in_bits[15:8] : _GEN_44; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_189 = 8'h2c == _T_4 ? io_in_bits[15:8] : _GEN_45; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_190 = 8'h2d == _T_4 ? io_in_bits[15:8] : _GEN_46; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_191 = 8'h2e == _T_4 ? io_in_bits[15:8] : _GEN_47; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_192 = 8'h2f == _T_4 ? io_in_bits[15:8] : _GEN_48; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_193 = 8'h30 == _T_4 ? io_in_bits[15:8] : _GEN_49; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_194 = 8'h31 == _T_4 ? io_in_bits[15:8] : _GEN_50; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_195 = 8'h32 == _T_4 ? io_in_bits[15:8] : _GEN_51; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_196 = 8'h33 == _T_4 ? io_in_bits[15:8] : _GEN_52; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_197 = 8'h34 == _T_4 ? io_in_bits[15:8] : _GEN_53; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_198 = 8'h35 == _T_4 ? io_in_bits[15:8] : _GEN_54; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_199 = 8'h36 == _T_4 ? io_in_bits[15:8] : _GEN_55; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_200 = 8'h37 == _T_4 ? io_in_bits[15:8] : _GEN_56; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_201 = 8'h38 == _T_4 ? io_in_bits[15:8] : _GEN_57; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_202 = 8'h39 == _T_4 ? io_in_bits[15:8] : _GEN_58; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_203 = 8'h3a == _T_4 ? io_in_bits[15:8] : _GEN_59; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_204 = 8'h3b == _T_4 ? io_in_bits[15:8] : _GEN_60; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_205 = 8'h3c == _T_4 ? io_in_bits[15:8] : _GEN_61; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_206 = 8'h3d == _T_4 ? io_in_bits[15:8] : _GEN_62; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_207 = 8'h3e == _T_4 ? io_in_bits[15:8] : _GEN_63; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_208 = 8'h3f == _T_4 ? io_in_bits[15:8] : _GEN_64; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_209 = 8'h40 == _T_4 ? io_in_bits[15:8] : _GEN_65; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_210 = 8'h41 == _T_4 ? io_in_bits[15:8] : _GEN_66; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_211 = 8'h42 == _T_4 ? io_in_bits[15:8] : _GEN_67; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_212 = 8'h43 == _T_4 ? io_in_bits[15:8] : _GEN_68; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_213 = 8'h44 == _T_4 ? io_in_bits[15:8] : _GEN_69; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_214 = 8'h45 == _T_4 ? io_in_bits[15:8] : _GEN_70; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_215 = 8'h46 == _T_4 ? io_in_bits[15:8] : _GEN_71; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_216 = 8'h47 == _T_4 ? io_in_bits[15:8] : _GEN_72; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_217 = 8'h48 == _T_4 ? io_in_bits[15:8] : _GEN_73; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_218 = 8'h49 == _T_4 ? io_in_bits[15:8] : _GEN_74; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_219 = 8'h4a == _T_4 ? io_in_bits[15:8] : _GEN_75; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_220 = 8'h4b == _T_4 ? io_in_bits[15:8] : _GEN_76; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_221 = 8'h4c == _T_4 ? io_in_bits[15:8] : _GEN_77; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_222 = 8'h4d == _T_4 ? io_in_bits[15:8] : _GEN_78; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_223 = 8'h4e == _T_4 ? io_in_bits[15:8] : _GEN_79; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_224 = 8'h4f == _T_4 ? io_in_bits[15:8] : _GEN_80; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_225 = 8'h50 == _T_4 ? io_in_bits[15:8] : _GEN_81; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_226 = 8'h51 == _T_4 ? io_in_bits[15:8] : _GEN_82; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_227 = 8'h52 == _T_4 ? io_in_bits[15:8] : _GEN_83; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_228 = 8'h53 == _T_4 ? io_in_bits[15:8] : _GEN_84; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_229 = 8'h54 == _T_4 ? io_in_bits[15:8] : _GEN_85; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_230 = 8'h55 == _T_4 ? io_in_bits[15:8] : _GEN_86; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_231 = 8'h56 == _T_4 ? io_in_bits[15:8] : _GEN_87; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_232 = 8'h57 == _T_4 ? io_in_bits[15:8] : _GEN_88; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_233 = 8'h58 == _T_4 ? io_in_bits[15:8] : _GEN_89; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_234 = 8'h59 == _T_4 ? io_in_bits[15:8] : _GEN_90; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_235 = 8'h5a == _T_4 ? io_in_bits[15:8] : _GEN_91; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_236 = 8'h5b == _T_4 ? io_in_bits[15:8] : _GEN_92; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_237 = 8'h5c == _T_4 ? io_in_bits[15:8] : _GEN_93; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_238 = 8'h5d == _T_4 ? io_in_bits[15:8] : _GEN_94; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_239 = 8'h5e == _T_4 ? io_in_bits[15:8] : _GEN_95; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_240 = 8'h5f == _T_4 ? io_in_bits[15:8] : _GEN_96; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_241 = 8'h60 == _T_4 ? io_in_bits[15:8] : _GEN_97; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_242 = 8'h61 == _T_4 ? io_in_bits[15:8] : _GEN_98; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_243 = 8'h62 == _T_4 ? io_in_bits[15:8] : _GEN_99; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_244 = 8'h63 == _T_4 ? io_in_bits[15:8] : _GEN_100; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_245 = 8'h64 == _T_4 ? io_in_bits[15:8] : _GEN_101; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_246 = 8'h65 == _T_4 ? io_in_bits[15:8] : _GEN_102; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_247 = 8'h66 == _T_4 ? io_in_bits[15:8] : _GEN_103; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_248 = 8'h67 == _T_4 ? io_in_bits[15:8] : _GEN_104; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_249 = 8'h68 == _T_4 ? io_in_bits[15:8] : _GEN_105; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_250 = 8'h69 == _T_4 ? io_in_bits[15:8] : _GEN_106; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_251 = 8'h6a == _T_4 ? io_in_bits[15:8] : _GEN_107; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_252 = 8'h6b == _T_4 ? io_in_bits[15:8] : _GEN_108; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_253 = 8'h6c == _T_4 ? io_in_bits[15:8] : _GEN_109; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_254 = 8'h6d == _T_4 ? io_in_bits[15:8] : _GEN_110; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_255 = 8'h6e == _T_4 ? io_in_bits[15:8] : _GEN_111; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_256 = 8'h6f == _T_4 ? io_in_bits[15:8] : _GEN_112; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_257 = 8'h70 == _T_4 ? io_in_bits[15:8] : _GEN_113; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_258 = 8'h71 == _T_4 ? io_in_bits[15:8] : _GEN_114; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_259 = 8'h72 == _T_4 ? io_in_bits[15:8] : _GEN_115; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_260 = 8'h73 == _T_4 ? io_in_bits[15:8] : _GEN_116; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_261 = 8'h74 == _T_4 ? io_in_bits[15:8] : _GEN_117; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_262 = 8'h75 == _T_4 ? io_in_bits[15:8] : _GEN_118; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_263 = 8'h76 == _T_4 ? io_in_bits[15:8] : _GEN_119; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_264 = 8'h77 == _T_4 ? io_in_bits[15:8] : _GEN_120; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_265 = 8'h78 == _T_4 ? io_in_bits[15:8] : _GEN_121; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_266 = 8'h79 == _T_4 ? io_in_bits[15:8] : _GEN_122; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_267 = 8'h7a == _T_4 ? io_in_bits[15:8] : _GEN_123; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_268 = 8'h7b == _T_4 ? io_in_bits[15:8] : _GEN_124; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_269 = 8'h7c == _T_4 ? io_in_bits[15:8] : _GEN_125; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_270 = 8'h7d == _T_4 ? io_in_bits[15:8] : _GEN_126; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_271 = 8'h7e == _T_4 ? io_in_bits[15:8] : _GEN_127; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_272 = 8'h7f == _T_4 ? io_in_bits[15:8] : _GEN_128; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_273 = 8'h80 == _T_4 ? io_in_bits[15:8] : _GEN_129; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_274 = 8'h81 == _T_4 ? io_in_bits[15:8] : _GEN_130; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_275 = 8'h82 == _T_4 ? io_in_bits[15:8] : _GEN_131; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_276 = 8'h83 == _T_4 ? io_in_bits[15:8] : _GEN_132; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_277 = 8'h84 == _T_4 ? io_in_bits[15:8] : _GEN_133; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_278 = 8'h85 == _T_4 ? io_in_bits[15:8] : _GEN_134; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_279 = 8'h86 == _T_4 ? io_in_bits[15:8] : _GEN_135; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_280 = 8'h87 == _T_4 ? io_in_bits[15:8] : _GEN_136; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_281 = 8'h88 == _T_4 ? io_in_bits[15:8] : _GEN_137; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_282 = 8'h89 == _T_4 ? io_in_bits[15:8] : _GEN_138; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_283 = 8'h8a == _T_4 ? io_in_bits[15:8] : _GEN_139; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_284 = 8'h8b == _T_4 ? io_in_bits[15:8] : _GEN_140; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_285 = 8'h8c == _T_4 ? io_in_bits[15:8] : _GEN_141; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_286 = 8'h8d == _T_4 ? io_in_bits[15:8] : _GEN_142; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_287 = 8'h8e == _T_4 ? io_in_bits[15:8] : _GEN_143; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_288 = 8'h8f == _T_4 ? io_in_bits[15:8] : _GEN_144; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_6 = enqPtr + 8'h2; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_289 = 8'h0 == _T_6 ? io_in_bits[23:16] : _GEN_145; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_290 = 8'h1 == _T_6 ? io_in_bits[23:16] : _GEN_146; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_291 = 8'h2 == _T_6 ? io_in_bits[23:16] : _GEN_147; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_292 = 8'h3 == _T_6 ? io_in_bits[23:16] : _GEN_148; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_293 = 8'h4 == _T_6 ? io_in_bits[23:16] : _GEN_149; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_294 = 8'h5 == _T_6 ? io_in_bits[23:16] : _GEN_150; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_295 = 8'h6 == _T_6 ? io_in_bits[23:16] : _GEN_151; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_296 = 8'h7 == _T_6 ? io_in_bits[23:16] : _GEN_152; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_297 = 8'h8 == _T_6 ? io_in_bits[23:16] : _GEN_153; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_298 = 8'h9 == _T_6 ? io_in_bits[23:16] : _GEN_154; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_299 = 8'ha == _T_6 ? io_in_bits[23:16] : _GEN_155; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_300 = 8'hb == _T_6 ? io_in_bits[23:16] : _GEN_156; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_301 = 8'hc == _T_6 ? io_in_bits[23:16] : _GEN_157; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_302 = 8'hd == _T_6 ? io_in_bits[23:16] : _GEN_158; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_303 = 8'he == _T_6 ? io_in_bits[23:16] : _GEN_159; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_304 = 8'hf == _T_6 ? io_in_bits[23:16] : _GEN_160; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_305 = 8'h10 == _T_6 ? io_in_bits[23:16] : _GEN_161; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_306 = 8'h11 == _T_6 ? io_in_bits[23:16] : _GEN_162; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_307 = 8'h12 == _T_6 ? io_in_bits[23:16] : _GEN_163; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_308 = 8'h13 == _T_6 ? io_in_bits[23:16] : _GEN_164; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_309 = 8'h14 == _T_6 ? io_in_bits[23:16] : _GEN_165; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_310 = 8'h15 == _T_6 ? io_in_bits[23:16] : _GEN_166; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_311 = 8'h16 == _T_6 ? io_in_bits[23:16] : _GEN_167; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_312 = 8'h17 == _T_6 ? io_in_bits[23:16] : _GEN_168; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_313 = 8'h18 == _T_6 ? io_in_bits[23:16] : _GEN_169; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_314 = 8'h19 == _T_6 ? io_in_bits[23:16] : _GEN_170; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_315 = 8'h1a == _T_6 ? io_in_bits[23:16] : _GEN_171; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_316 = 8'h1b == _T_6 ? io_in_bits[23:16] : _GEN_172; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_317 = 8'h1c == _T_6 ? io_in_bits[23:16] : _GEN_173; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_318 = 8'h1d == _T_6 ? io_in_bits[23:16] : _GEN_174; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_319 = 8'h1e == _T_6 ? io_in_bits[23:16] : _GEN_175; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_320 = 8'h1f == _T_6 ? io_in_bits[23:16] : _GEN_176; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_321 = 8'h20 == _T_6 ? io_in_bits[23:16] : _GEN_177; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_322 = 8'h21 == _T_6 ? io_in_bits[23:16] : _GEN_178; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_323 = 8'h22 == _T_6 ? io_in_bits[23:16] : _GEN_179; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_324 = 8'h23 == _T_6 ? io_in_bits[23:16] : _GEN_180; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_325 = 8'h24 == _T_6 ? io_in_bits[23:16] : _GEN_181; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_326 = 8'h25 == _T_6 ? io_in_bits[23:16] : _GEN_182; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_327 = 8'h26 == _T_6 ? io_in_bits[23:16] : _GEN_183; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_328 = 8'h27 == _T_6 ? io_in_bits[23:16] : _GEN_184; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_329 = 8'h28 == _T_6 ? io_in_bits[23:16] : _GEN_185; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_330 = 8'h29 == _T_6 ? io_in_bits[23:16] : _GEN_186; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_331 = 8'h2a == _T_6 ? io_in_bits[23:16] : _GEN_187; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_332 = 8'h2b == _T_6 ? io_in_bits[23:16] : _GEN_188; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_333 = 8'h2c == _T_6 ? io_in_bits[23:16] : _GEN_189; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_334 = 8'h2d == _T_6 ? io_in_bits[23:16] : _GEN_190; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_335 = 8'h2e == _T_6 ? io_in_bits[23:16] : _GEN_191; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_336 = 8'h2f == _T_6 ? io_in_bits[23:16] : _GEN_192; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_337 = 8'h30 == _T_6 ? io_in_bits[23:16] : _GEN_193; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_338 = 8'h31 == _T_6 ? io_in_bits[23:16] : _GEN_194; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_339 = 8'h32 == _T_6 ? io_in_bits[23:16] : _GEN_195; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_340 = 8'h33 == _T_6 ? io_in_bits[23:16] : _GEN_196; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_341 = 8'h34 == _T_6 ? io_in_bits[23:16] : _GEN_197; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_342 = 8'h35 == _T_6 ? io_in_bits[23:16] : _GEN_198; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_343 = 8'h36 == _T_6 ? io_in_bits[23:16] : _GEN_199; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_344 = 8'h37 == _T_6 ? io_in_bits[23:16] : _GEN_200; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_345 = 8'h38 == _T_6 ? io_in_bits[23:16] : _GEN_201; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_346 = 8'h39 == _T_6 ? io_in_bits[23:16] : _GEN_202; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_347 = 8'h3a == _T_6 ? io_in_bits[23:16] : _GEN_203; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_348 = 8'h3b == _T_6 ? io_in_bits[23:16] : _GEN_204; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_349 = 8'h3c == _T_6 ? io_in_bits[23:16] : _GEN_205; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_350 = 8'h3d == _T_6 ? io_in_bits[23:16] : _GEN_206; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_351 = 8'h3e == _T_6 ? io_in_bits[23:16] : _GEN_207; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_352 = 8'h3f == _T_6 ? io_in_bits[23:16] : _GEN_208; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_353 = 8'h40 == _T_6 ? io_in_bits[23:16] : _GEN_209; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_354 = 8'h41 == _T_6 ? io_in_bits[23:16] : _GEN_210; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_355 = 8'h42 == _T_6 ? io_in_bits[23:16] : _GEN_211; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_356 = 8'h43 == _T_6 ? io_in_bits[23:16] : _GEN_212; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_357 = 8'h44 == _T_6 ? io_in_bits[23:16] : _GEN_213; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_358 = 8'h45 == _T_6 ? io_in_bits[23:16] : _GEN_214; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_359 = 8'h46 == _T_6 ? io_in_bits[23:16] : _GEN_215; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_360 = 8'h47 == _T_6 ? io_in_bits[23:16] : _GEN_216; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_361 = 8'h48 == _T_6 ? io_in_bits[23:16] : _GEN_217; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_362 = 8'h49 == _T_6 ? io_in_bits[23:16] : _GEN_218; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_363 = 8'h4a == _T_6 ? io_in_bits[23:16] : _GEN_219; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_364 = 8'h4b == _T_6 ? io_in_bits[23:16] : _GEN_220; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_365 = 8'h4c == _T_6 ? io_in_bits[23:16] : _GEN_221; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_366 = 8'h4d == _T_6 ? io_in_bits[23:16] : _GEN_222; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_367 = 8'h4e == _T_6 ? io_in_bits[23:16] : _GEN_223; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_368 = 8'h4f == _T_6 ? io_in_bits[23:16] : _GEN_224; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_369 = 8'h50 == _T_6 ? io_in_bits[23:16] : _GEN_225; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_370 = 8'h51 == _T_6 ? io_in_bits[23:16] : _GEN_226; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_371 = 8'h52 == _T_6 ? io_in_bits[23:16] : _GEN_227; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_372 = 8'h53 == _T_6 ? io_in_bits[23:16] : _GEN_228; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_373 = 8'h54 == _T_6 ? io_in_bits[23:16] : _GEN_229; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_374 = 8'h55 == _T_6 ? io_in_bits[23:16] : _GEN_230; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_375 = 8'h56 == _T_6 ? io_in_bits[23:16] : _GEN_231; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_376 = 8'h57 == _T_6 ? io_in_bits[23:16] : _GEN_232; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_377 = 8'h58 == _T_6 ? io_in_bits[23:16] : _GEN_233; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_378 = 8'h59 == _T_6 ? io_in_bits[23:16] : _GEN_234; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_379 = 8'h5a == _T_6 ? io_in_bits[23:16] : _GEN_235; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_380 = 8'h5b == _T_6 ? io_in_bits[23:16] : _GEN_236; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_381 = 8'h5c == _T_6 ? io_in_bits[23:16] : _GEN_237; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_382 = 8'h5d == _T_6 ? io_in_bits[23:16] : _GEN_238; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_383 = 8'h5e == _T_6 ? io_in_bits[23:16] : _GEN_239; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_384 = 8'h5f == _T_6 ? io_in_bits[23:16] : _GEN_240; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_385 = 8'h60 == _T_6 ? io_in_bits[23:16] : _GEN_241; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_386 = 8'h61 == _T_6 ? io_in_bits[23:16] : _GEN_242; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_387 = 8'h62 == _T_6 ? io_in_bits[23:16] : _GEN_243; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_388 = 8'h63 == _T_6 ? io_in_bits[23:16] : _GEN_244; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_389 = 8'h64 == _T_6 ? io_in_bits[23:16] : _GEN_245; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_390 = 8'h65 == _T_6 ? io_in_bits[23:16] : _GEN_246; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_391 = 8'h66 == _T_6 ? io_in_bits[23:16] : _GEN_247; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_392 = 8'h67 == _T_6 ? io_in_bits[23:16] : _GEN_248; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_393 = 8'h68 == _T_6 ? io_in_bits[23:16] : _GEN_249; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_394 = 8'h69 == _T_6 ? io_in_bits[23:16] : _GEN_250; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_395 = 8'h6a == _T_6 ? io_in_bits[23:16] : _GEN_251; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_396 = 8'h6b == _T_6 ? io_in_bits[23:16] : _GEN_252; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_397 = 8'h6c == _T_6 ? io_in_bits[23:16] : _GEN_253; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_398 = 8'h6d == _T_6 ? io_in_bits[23:16] : _GEN_254; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_399 = 8'h6e == _T_6 ? io_in_bits[23:16] : _GEN_255; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_400 = 8'h6f == _T_6 ? io_in_bits[23:16] : _GEN_256; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_401 = 8'h70 == _T_6 ? io_in_bits[23:16] : _GEN_257; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_402 = 8'h71 == _T_6 ? io_in_bits[23:16] : _GEN_258; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_403 = 8'h72 == _T_6 ? io_in_bits[23:16] : _GEN_259; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_404 = 8'h73 == _T_6 ? io_in_bits[23:16] : _GEN_260; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_405 = 8'h74 == _T_6 ? io_in_bits[23:16] : _GEN_261; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_406 = 8'h75 == _T_6 ? io_in_bits[23:16] : _GEN_262; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_407 = 8'h76 == _T_6 ? io_in_bits[23:16] : _GEN_263; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_408 = 8'h77 == _T_6 ? io_in_bits[23:16] : _GEN_264; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_409 = 8'h78 == _T_6 ? io_in_bits[23:16] : _GEN_265; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_410 = 8'h79 == _T_6 ? io_in_bits[23:16] : _GEN_266; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_411 = 8'h7a == _T_6 ? io_in_bits[23:16] : _GEN_267; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_412 = 8'h7b == _T_6 ? io_in_bits[23:16] : _GEN_268; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_413 = 8'h7c == _T_6 ? io_in_bits[23:16] : _GEN_269; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_414 = 8'h7d == _T_6 ? io_in_bits[23:16] : _GEN_270; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_415 = 8'h7e == _T_6 ? io_in_bits[23:16] : _GEN_271; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_416 = 8'h7f == _T_6 ? io_in_bits[23:16] : _GEN_272; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_417 = 8'h80 == _T_6 ? io_in_bits[23:16] : _GEN_273; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_418 = 8'h81 == _T_6 ? io_in_bits[23:16] : _GEN_274; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_419 = 8'h82 == _T_6 ? io_in_bits[23:16] : _GEN_275; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_420 = 8'h83 == _T_6 ? io_in_bits[23:16] : _GEN_276; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_421 = 8'h84 == _T_6 ? io_in_bits[23:16] : _GEN_277; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_422 = 8'h85 == _T_6 ? io_in_bits[23:16] : _GEN_278; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_423 = 8'h86 == _T_6 ? io_in_bits[23:16] : _GEN_279; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_424 = 8'h87 == _T_6 ? io_in_bits[23:16] : _GEN_280; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_425 = 8'h88 == _T_6 ? io_in_bits[23:16] : _GEN_281; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_426 = 8'h89 == _T_6 ? io_in_bits[23:16] : _GEN_282; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_427 = 8'h8a == _T_6 ? io_in_bits[23:16] : _GEN_283; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_428 = 8'h8b == _T_6 ? io_in_bits[23:16] : _GEN_284; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_429 = 8'h8c == _T_6 ? io_in_bits[23:16] : _GEN_285; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_430 = 8'h8d == _T_6 ? io_in_bits[23:16] : _GEN_286; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_431 = 8'h8e == _T_6 ? io_in_bits[23:16] : _GEN_287; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_432 = 8'h8f == _T_6 ? io_in_bits[23:16] : _GEN_288; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_8 = enqPtr + 8'h3; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_433 = 8'h0 == _T_8 ? io_in_bits[31:24] : _GEN_289; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_434 = 8'h1 == _T_8 ? io_in_bits[31:24] : _GEN_290; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_435 = 8'h2 == _T_8 ? io_in_bits[31:24] : _GEN_291; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_436 = 8'h3 == _T_8 ? io_in_bits[31:24] : _GEN_292; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_437 = 8'h4 == _T_8 ? io_in_bits[31:24] : _GEN_293; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_438 = 8'h5 == _T_8 ? io_in_bits[31:24] : _GEN_294; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_439 = 8'h6 == _T_8 ? io_in_bits[31:24] : _GEN_295; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_440 = 8'h7 == _T_8 ? io_in_bits[31:24] : _GEN_296; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_441 = 8'h8 == _T_8 ? io_in_bits[31:24] : _GEN_297; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_442 = 8'h9 == _T_8 ? io_in_bits[31:24] : _GEN_298; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_443 = 8'ha == _T_8 ? io_in_bits[31:24] : _GEN_299; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_444 = 8'hb == _T_8 ? io_in_bits[31:24] : _GEN_300; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_445 = 8'hc == _T_8 ? io_in_bits[31:24] : _GEN_301; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_446 = 8'hd == _T_8 ? io_in_bits[31:24] : _GEN_302; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_447 = 8'he == _T_8 ? io_in_bits[31:24] : _GEN_303; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_448 = 8'hf == _T_8 ? io_in_bits[31:24] : _GEN_304; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_449 = 8'h10 == _T_8 ? io_in_bits[31:24] : _GEN_305; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_450 = 8'h11 == _T_8 ? io_in_bits[31:24] : _GEN_306; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_451 = 8'h12 == _T_8 ? io_in_bits[31:24] : _GEN_307; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_452 = 8'h13 == _T_8 ? io_in_bits[31:24] : _GEN_308; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_453 = 8'h14 == _T_8 ? io_in_bits[31:24] : _GEN_309; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_454 = 8'h15 == _T_8 ? io_in_bits[31:24] : _GEN_310; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_455 = 8'h16 == _T_8 ? io_in_bits[31:24] : _GEN_311; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_456 = 8'h17 == _T_8 ? io_in_bits[31:24] : _GEN_312; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_457 = 8'h18 == _T_8 ? io_in_bits[31:24] : _GEN_313; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_458 = 8'h19 == _T_8 ? io_in_bits[31:24] : _GEN_314; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_459 = 8'h1a == _T_8 ? io_in_bits[31:24] : _GEN_315; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_460 = 8'h1b == _T_8 ? io_in_bits[31:24] : _GEN_316; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_461 = 8'h1c == _T_8 ? io_in_bits[31:24] : _GEN_317; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_462 = 8'h1d == _T_8 ? io_in_bits[31:24] : _GEN_318; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_463 = 8'h1e == _T_8 ? io_in_bits[31:24] : _GEN_319; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_464 = 8'h1f == _T_8 ? io_in_bits[31:24] : _GEN_320; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_465 = 8'h20 == _T_8 ? io_in_bits[31:24] : _GEN_321; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_466 = 8'h21 == _T_8 ? io_in_bits[31:24] : _GEN_322; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_467 = 8'h22 == _T_8 ? io_in_bits[31:24] : _GEN_323; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_468 = 8'h23 == _T_8 ? io_in_bits[31:24] : _GEN_324; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_469 = 8'h24 == _T_8 ? io_in_bits[31:24] : _GEN_325; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_470 = 8'h25 == _T_8 ? io_in_bits[31:24] : _GEN_326; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_471 = 8'h26 == _T_8 ? io_in_bits[31:24] : _GEN_327; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_472 = 8'h27 == _T_8 ? io_in_bits[31:24] : _GEN_328; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_473 = 8'h28 == _T_8 ? io_in_bits[31:24] : _GEN_329; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_474 = 8'h29 == _T_8 ? io_in_bits[31:24] : _GEN_330; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_475 = 8'h2a == _T_8 ? io_in_bits[31:24] : _GEN_331; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_476 = 8'h2b == _T_8 ? io_in_bits[31:24] : _GEN_332; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_477 = 8'h2c == _T_8 ? io_in_bits[31:24] : _GEN_333; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_478 = 8'h2d == _T_8 ? io_in_bits[31:24] : _GEN_334; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_479 = 8'h2e == _T_8 ? io_in_bits[31:24] : _GEN_335; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_480 = 8'h2f == _T_8 ? io_in_bits[31:24] : _GEN_336; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_481 = 8'h30 == _T_8 ? io_in_bits[31:24] : _GEN_337; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_482 = 8'h31 == _T_8 ? io_in_bits[31:24] : _GEN_338; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_483 = 8'h32 == _T_8 ? io_in_bits[31:24] : _GEN_339; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_484 = 8'h33 == _T_8 ? io_in_bits[31:24] : _GEN_340; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_485 = 8'h34 == _T_8 ? io_in_bits[31:24] : _GEN_341; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_486 = 8'h35 == _T_8 ? io_in_bits[31:24] : _GEN_342; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_487 = 8'h36 == _T_8 ? io_in_bits[31:24] : _GEN_343; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_488 = 8'h37 == _T_8 ? io_in_bits[31:24] : _GEN_344; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_489 = 8'h38 == _T_8 ? io_in_bits[31:24] : _GEN_345; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_490 = 8'h39 == _T_8 ? io_in_bits[31:24] : _GEN_346; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_491 = 8'h3a == _T_8 ? io_in_bits[31:24] : _GEN_347; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_492 = 8'h3b == _T_8 ? io_in_bits[31:24] : _GEN_348; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_493 = 8'h3c == _T_8 ? io_in_bits[31:24] : _GEN_349; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_494 = 8'h3d == _T_8 ? io_in_bits[31:24] : _GEN_350; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_495 = 8'h3e == _T_8 ? io_in_bits[31:24] : _GEN_351; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_496 = 8'h3f == _T_8 ? io_in_bits[31:24] : _GEN_352; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_497 = 8'h40 == _T_8 ? io_in_bits[31:24] : _GEN_353; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_498 = 8'h41 == _T_8 ? io_in_bits[31:24] : _GEN_354; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_499 = 8'h42 == _T_8 ? io_in_bits[31:24] : _GEN_355; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_500 = 8'h43 == _T_8 ? io_in_bits[31:24] : _GEN_356; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_501 = 8'h44 == _T_8 ? io_in_bits[31:24] : _GEN_357; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_502 = 8'h45 == _T_8 ? io_in_bits[31:24] : _GEN_358; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_503 = 8'h46 == _T_8 ? io_in_bits[31:24] : _GEN_359; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_504 = 8'h47 == _T_8 ? io_in_bits[31:24] : _GEN_360; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_505 = 8'h48 == _T_8 ? io_in_bits[31:24] : _GEN_361; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_506 = 8'h49 == _T_8 ? io_in_bits[31:24] : _GEN_362; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_507 = 8'h4a == _T_8 ? io_in_bits[31:24] : _GEN_363; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_508 = 8'h4b == _T_8 ? io_in_bits[31:24] : _GEN_364; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_509 = 8'h4c == _T_8 ? io_in_bits[31:24] : _GEN_365; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_510 = 8'h4d == _T_8 ? io_in_bits[31:24] : _GEN_366; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_511 = 8'h4e == _T_8 ? io_in_bits[31:24] : _GEN_367; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_512 = 8'h4f == _T_8 ? io_in_bits[31:24] : _GEN_368; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_513 = 8'h50 == _T_8 ? io_in_bits[31:24] : _GEN_369; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_514 = 8'h51 == _T_8 ? io_in_bits[31:24] : _GEN_370; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_515 = 8'h52 == _T_8 ? io_in_bits[31:24] : _GEN_371; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_516 = 8'h53 == _T_8 ? io_in_bits[31:24] : _GEN_372; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_517 = 8'h54 == _T_8 ? io_in_bits[31:24] : _GEN_373; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_518 = 8'h55 == _T_8 ? io_in_bits[31:24] : _GEN_374; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_519 = 8'h56 == _T_8 ? io_in_bits[31:24] : _GEN_375; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_520 = 8'h57 == _T_8 ? io_in_bits[31:24] : _GEN_376; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_521 = 8'h58 == _T_8 ? io_in_bits[31:24] : _GEN_377; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_522 = 8'h59 == _T_8 ? io_in_bits[31:24] : _GEN_378; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_523 = 8'h5a == _T_8 ? io_in_bits[31:24] : _GEN_379; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_524 = 8'h5b == _T_8 ? io_in_bits[31:24] : _GEN_380; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_525 = 8'h5c == _T_8 ? io_in_bits[31:24] : _GEN_381; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_526 = 8'h5d == _T_8 ? io_in_bits[31:24] : _GEN_382; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_527 = 8'h5e == _T_8 ? io_in_bits[31:24] : _GEN_383; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_528 = 8'h5f == _T_8 ? io_in_bits[31:24] : _GEN_384; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_529 = 8'h60 == _T_8 ? io_in_bits[31:24] : _GEN_385; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_530 = 8'h61 == _T_8 ? io_in_bits[31:24] : _GEN_386; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_531 = 8'h62 == _T_8 ? io_in_bits[31:24] : _GEN_387; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_532 = 8'h63 == _T_8 ? io_in_bits[31:24] : _GEN_388; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_533 = 8'h64 == _T_8 ? io_in_bits[31:24] : _GEN_389; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_534 = 8'h65 == _T_8 ? io_in_bits[31:24] : _GEN_390; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_535 = 8'h66 == _T_8 ? io_in_bits[31:24] : _GEN_391; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_536 = 8'h67 == _T_8 ? io_in_bits[31:24] : _GEN_392; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_537 = 8'h68 == _T_8 ? io_in_bits[31:24] : _GEN_393; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_538 = 8'h69 == _T_8 ? io_in_bits[31:24] : _GEN_394; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_539 = 8'h6a == _T_8 ? io_in_bits[31:24] : _GEN_395; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_540 = 8'h6b == _T_8 ? io_in_bits[31:24] : _GEN_396; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_541 = 8'h6c == _T_8 ? io_in_bits[31:24] : _GEN_397; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_542 = 8'h6d == _T_8 ? io_in_bits[31:24] : _GEN_398; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_543 = 8'h6e == _T_8 ? io_in_bits[31:24] : _GEN_399; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_544 = 8'h6f == _T_8 ? io_in_bits[31:24] : _GEN_400; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_545 = 8'h70 == _T_8 ? io_in_bits[31:24] : _GEN_401; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_546 = 8'h71 == _T_8 ? io_in_bits[31:24] : _GEN_402; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_547 = 8'h72 == _T_8 ? io_in_bits[31:24] : _GEN_403; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_548 = 8'h73 == _T_8 ? io_in_bits[31:24] : _GEN_404; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_549 = 8'h74 == _T_8 ? io_in_bits[31:24] : _GEN_405; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_550 = 8'h75 == _T_8 ? io_in_bits[31:24] : _GEN_406; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_551 = 8'h76 == _T_8 ? io_in_bits[31:24] : _GEN_407; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_552 = 8'h77 == _T_8 ? io_in_bits[31:24] : _GEN_408; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_553 = 8'h78 == _T_8 ? io_in_bits[31:24] : _GEN_409; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_554 = 8'h79 == _T_8 ? io_in_bits[31:24] : _GEN_410; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_555 = 8'h7a == _T_8 ? io_in_bits[31:24] : _GEN_411; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_556 = 8'h7b == _T_8 ? io_in_bits[31:24] : _GEN_412; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_557 = 8'h7c == _T_8 ? io_in_bits[31:24] : _GEN_413; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_558 = 8'h7d == _T_8 ? io_in_bits[31:24] : _GEN_414; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_559 = 8'h7e == _T_8 ? io_in_bits[31:24] : _GEN_415; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_560 = 8'h7f == _T_8 ? io_in_bits[31:24] : _GEN_416; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_561 = 8'h80 == _T_8 ? io_in_bits[31:24] : _GEN_417; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_562 = 8'h81 == _T_8 ? io_in_bits[31:24] : _GEN_418; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_563 = 8'h82 == _T_8 ? io_in_bits[31:24] : _GEN_419; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_564 = 8'h83 == _T_8 ? io_in_bits[31:24] : _GEN_420; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_565 = 8'h84 == _T_8 ? io_in_bits[31:24] : _GEN_421; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_566 = 8'h85 == _T_8 ? io_in_bits[31:24] : _GEN_422; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_567 = 8'h86 == _T_8 ? io_in_bits[31:24] : _GEN_423; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_568 = 8'h87 == _T_8 ? io_in_bits[31:24] : _GEN_424; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_569 = 8'h88 == _T_8 ? io_in_bits[31:24] : _GEN_425; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_570 = 8'h89 == _T_8 ? io_in_bits[31:24] : _GEN_426; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_571 = 8'h8a == _T_8 ? io_in_bits[31:24] : _GEN_427; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_572 = 8'h8b == _T_8 ? io_in_bits[31:24] : _GEN_428; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_573 = 8'h8c == _T_8 ? io_in_bits[31:24] : _GEN_429; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_574 = 8'h8d == _T_8 ? io_in_bits[31:24] : _GEN_430; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_575 = 8'h8e == _T_8 ? io_in_bits[31:24] : _GEN_431; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_576 = 8'h8f == _T_8 ? io_in_bits[31:24] : _GEN_432; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_10 = enqPtr + 8'h4; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_577 = 8'h0 == _T_10 ? io_in_bits[39:32] : _GEN_433; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_578 = 8'h1 == _T_10 ? io_in_bits[39:32] : _GEN_434; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_579 = 8'h2 == _T_10 ? io_in_bits[39:32] : _GEN_435; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_580 = 8'h3 == _T_10 ? io_in_bits[39:32] : _GEN_436; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_581 = 8'h4 == _T_10 ? io_in_bits[39:32] : _GEN_437; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_582 = 8'h5 == _T_10 ? io_in_bits[39:32] : _GEN_438; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_583 = 8'h6 == _T_10 ? io_in_bits[39:32] : _GEN_439; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_584 = 8'h7 == _T_10 ? io_in_bits[39:32] : _GEN_440; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_585 = 8'h8 == _T_10 ? io_in_bits[39:32] : _GEN_441; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_586 = 8'h9 == _T_10 ? io_in_bits[39:32] : _GEN_442; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_587 = 8'ha == _T_10 ? io_in_bits[39:32] : _GEN_443; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_588 = 8'hb == _T_10 ? io_in_bits[39:32] : _GEN_444; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_589 = 8'hc == _T_10 ? io_in_bits[39:32] : _GEN_445; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_590 = 8'hd == _T_10 ? io_in_bits[39:32] : _GEN_446; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_591 = 8'he == _T_10 ? io_in_bits[39:32] : _GEN_447; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_592 = 8'hf == _T_10 ? io_in_bits[39:32] : _GEN_448; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_593 = 8'h10 == _T_10 ? io_in_bits[39:32] : _GEN_449; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_594 = 8'h11 == _T_10 ? io_in_bits[39:32] : _GEN_450; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_595 = 8'h12 == _T_10 ? io_in_bits[39:32] : _GEN_451; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_596 = 8'h13 == _T_10 ? io_in_bits[39:32] : _GEN_452; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_597 = 8'h14 == _T_10 ? io_in_bits[39:32] : _GEN_453; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_598 = 8'h15 == _T_10 ? io_in_bits[39:32] : _GEN_454; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_599 = 8'h16 == _T_10 ? io_in_bits[39:32] : _GEN_455; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_600 = 8'h17 == _T_10 ? io_in_bits[39:32] : _GEN_456; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_601 = 8'h18 == _T_10 ? io_in_bits[39:32] : _GEN_457; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_602 = 8'h19 == _T_10 ? io_in_bits[39:32] : _GEN_458; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_603 = 8'h1a == _T_10 ? io_in_bits[39:32] : _GEN_459; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_604 = 8'h1b == _T_10 ? io_in_bits[39:32] : _GEN_460; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_605 = 8'h1c == _T_10 ? io_in_bits[39:32] : _GEN_461; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_606 = 8'h1d == _T_10 ? io_in_bits[39:32] : _GEN_462; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_607 = 8'h1e == _T_10 ? io_in_bits[39:32] : _GEN_463; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_608 = 8'h1f == _T_10 ? io_in_bits[39:32] : _GEN_464; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_609 = 8'h20 == _T_10 ? io_in_bits[39:32] : _GEN_465; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_610 = 8'h21 == _T_10 ? io_in_bits[39:32] : _GEN_466; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_611 = 8'h22 == _T_10 ? io_in_bits[39:32] : _GEN_467; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_612 = 8'h23 == _T_10 ? io_in_bits[39:32] : _GEN_468; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_613 = 8'h24 == _T_10 ? io_in_bits[39:32] : _GEN_469; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_614 = 8'h25 == _T_10 ? io_in_bits[39:32] : _GEN_470; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_615 = 8'h26 == _T_10 ? io_in_bits[39:32] : _GEN_471; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_616 = 8'h27 == _T_10 ? io_in_bits[39:32] : _GEN_472; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_617 = 8'h28 == _T_10 ? io_in_bits[39:32] : _GEN_473; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_618 = 8'h29 == _T_10 ? io_in_bits[39:32] : _GEN_474; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_619 = 8'h2a == _T_10 ? io_in_bits[39:32] : _GEN_475; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_620 = 8'h2b == _T_10 ? io_in_bits[39:32] : _GEN_476; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_621 = 8'h2c == _T_10 ? io_in_bits[39:32] : _GEN_477; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_622 = 8'h2d == _T_10 ? io_in_bits[39:32] : _GEN_478; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_623 = 8'h2e == _T_10 ? io_in_bits[39:32] : _GEN_479; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_624 = 8'h2f == _T_10 ? io_in_bits[39:32] : _GEN_480; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_625 = 8'h30 == _T_10 ? io_in_bits[39:32] : _GEN_481; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_626 = 8'h31 == _T_10 ? io_in_bits[39:32] : _GEN_482; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_627 = 8'h32 == _T_10 ? io_in_bits[39:32] : _GEN_483; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_628 = 8'h33 == _T_10 ? io_in_bits[39:32] : _GEN_484; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_629 = 8'h34 == _T_10 ? io_in_bits[39:32] : _GEN_485; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_630 = 8'h35 == _T_10 ? io_in_bits[39:32] : _GEN_486; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_631 = 8'h36 == _T_10 ? io_in_bits[39:32] : _GEN_487; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_632 = 8'h37 == _T_10 ? io_in_bits[39:32] : _GEN_488; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_633 = 8'h38 == _T_10 ? io_in_bits[39:32] : _GEN_489; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_634 = 8'h39 == _T_10 ? io_in_bits[39:32] : _GEN_490; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_635 = 8'h3a == _T_10 ? io_in_bits[39:32] : _GEN_491; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_636 = 8'h3b == _T_10 ? io_in_bits[39:32] : _GEN_492; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_637 = 8'h3c == _T_10 ? io_in_bits[39:32] : _GEN_493; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_638 = 8'h3d == _T_10 ? io_in_bits[39:32] : _GEN_494; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_639 = 8'h3e == _T_10 ? io_in_bits[39:32] : _GEN_495; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_640 = 8'h3f == _T_10 ? io_in_bits[39:32] : _GEN_496; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_641 = 8'h40 == _T_10 ? io_in_bits[39:32] : _GEN_497; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_642 = 8'h41 == _T_10 ? io_in_bits[39:32] : _GEN_498; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_643 = 8'h42 == _T_10 ? io_in_bits[39:32] : _GEN_499; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_644 = 8'h43 == _T_10 ? io_in_bits[39:32] : _GEN_500; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_645 = 8'h44 == _T_10 ? io_in_bits[39:32] : _GEN_501; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_646 = 8'h45 == _T_10 ? io_in_bits[39:32] : _GEN_502; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_647 = 8'h46 == _T_10 ? io_in_bits[39:32] : _GEN_503; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_648 = 8'h47 == _T_10 ? io_in_bits[39:32] : _GEN_504; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_649 = 8'h48 == _T_10 ? io_in_bits[39:32] : _GEN_505; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_650 = 8'h49 == _T_10 ? io_in_bits[39:32] : _GEN_506; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_651 = 8'h4a == _T_10 ? io_in_bits[39:32] : _GEN_507; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_652 = 8'h4b == _T_10 ? io_in_bits[39:32] : _GEN_508; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_653 = 8'h4c == _T_10 ? io_in_bits[39:32] : _GEN_509; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_654 = 8'h4d == _T_10 ? io_in_bits[39:32] : _GEN_510; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_655 = 8'h4e == _T_10 ? io_in_bits[39:32] : _GEN_511; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_656 = 8'h4f == _T_10 ? io_in_bits[39:32] : _GEN_512; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_657 = 8'h50 == _T_10 ? io_in_bits[39:32] : _GEN_513; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_658 = 8'h51 == _T_10 ? io_in_bits[39:32] : _GEN_514; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_659 = 8'h52 == _T_10 ? io_in_bits[39:32] : _GEN_515; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_660 = 8'h53 == _T_10 ? io_in_bits[39:32] : _GEN_516; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_661 = 8'h54 == _T_10 ? io_in_bits[39:32] : _GEN_517; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_662 = 8'h55 == _T_10 ? io_in_bits[39:32] : _GEN_518; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_663 = 8'h56 == _T_10 ? io_in_bits[39:32] : _GEN_519; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_664 = 8'h57 == _T_10 ? io_in_bits[39:32] : _GEN_520; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_665 = 8'h58 == _T_10 ? io_in_bits[39:32] : _GEN_521; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_666 = 8'h59 == _T_10 ? io_in_bits[39:32] : _GEN_522; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_667 = 8'h5a == _T_10 ? io_in_bits[39:32] : _GEN_523; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_668 = 8'h5b == _T_10 ? io_in_bits[39:32] : _GEN_524; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_669 = 8'h5c == _T_10 ? io_in_bits[39:32] : _GEN_525; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_670 = 8'h5d == _T_10 ? io_in_bits[39:32] : _GEN_526; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_671 = 8'h5e == _T_10 ? io_in_bits[39:32] : _GEN_527; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_672 = 8'h5f == _T_10 ? io_in_bits[39:32] : _GEN_528; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_673 = 8'h60 == _T_10 ? io_in_bits[39:32] : _GEN_529; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_674 = 8'h61 == _T_10 ? io_in_bits[39:32] : _GEN_530; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_675 = 8'h62 == _T_10 ? io_in_bits[39:32] : _GEN_531; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_676 = 8'h63 == _T_10 ? io_in_bits[39:32] : _GEN_532; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_677 = 8'h64 == _T_10 ? io_in_bits[39:32] : _GEN_533; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_678 = 8'h65 == _T_10 ? io_in_bits[39:32] : _GEN_534; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_679 = 8'h66 == _T_10 ? io_in_bits[39:32] : _GEN_535; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_680 = 8'h67 == _T_10 ? io_in_bits[39:32] : _GEN_536; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_681 = 8'h68 == _T_10 ? io_in_bits[39:32] : _GEN_537; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_682 = 8'h69 == _T_10 ? io_in_bits[39:32] : _GEN_538; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_683 = 8'h6a == _T_10 ? io_in_bits[39:32] : _GEN_539; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_684 = 8'h6b == _T_10 ? io_in_bits[39:32] : _GEN_540; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_685 = 8'h6c == _T_10 ? io_in_bits[39:32] : _GEN_541; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_686 = 8'h6d == _T_10 ? io_in_bits[39:32] : _GEN_542; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_687 = 8'h6e == _T_10 ? io_in_bits[39:32] : _GEN_543; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_688 = 8'h6f == _T_10 ? io_in_bits[39:32] : _GEN_544; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_689 = 8'h70 == _T_10 ? io_in_bits[39:32] : _GEN_545; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_690 = 8'h71 == _T_10 ? io_in_bits[39:32] : _GEN_546; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_691 = 8'h72 == _T_10 ? io_in_bits[39:32] : _GEN_547; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_692 = 8'h73 == _T_10 ? io_in_bits[39:32] : _GEN_548; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_693 = 8'h74 == _T_10 ? io_in_bits[39:32] : _GEN_549; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_694 = 8'h75 == _T_10 ? io_in_bits[39:32] : _GEN_550; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_695 = 8'h76 == _T_10 ? io_in_bits[39:32] : _GEN_551; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_696 = 8'h77 == _T_10 ? io_in_bits[39:32] : _GEN_552; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_697 = 8'h78 == _T_10 ? io_in_bits[39:32] : _GEN_553; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_698 = 8'h79 == _T_10 ? io_in_bits[39:32] : _GEN_554; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_699 = 8'h7a == _T_10 ? io_in_bits[39:32] : _GEN_555; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_700 = 8'h7b == _T_10 ? io_in_bits[39:32] : _GEN_556; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_701 = 8'h7c == _T_10 ? io_in_bits[39:32] : _GEN_557; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_702 = 8'h7d == _T_10 ? io_in_bits[39:32] : _GEN_558; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_703 = 8'h7e == _T_10 ? io_in_bits[39:32] : _GEN_559; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_704 = 8'h7f == _T_10 ? io_in_bits[39:32] : _GEN_560; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_705 = 8'h80 == _T_10 ? io_in_bits[39:32] : _GEN_561; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_706 = 8'h81 == _T_10 ? io_in_bits[39:32] : _GEN_562; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_707 = 8'h82 == _T_10 ? io_in_bits[39:32] : _GEN_563; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_708 = 8'h83 == _T_10 ? io_in_bits[39:32] : _GEN_564; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_709 = 8'h84 == _T_10 ? io_in_bits[39:32] : _GEN_565; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_710 = 8'h85 == _T_10 ? io_in_bits[39:32] : _GEN_566; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_711 = 8'h86 == _T_10 ? io_in_bits[39:32] : _GEN_567; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_712 = 8'h87 == _T_10 ? io_in_bits[39:32] : _GEN_568; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_713 = 8'h88 == _T_10 ? io_in_bits[39:32] : _GEN_569; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_714 = 8'h89 == _T_10 ? io_in_bits[39:32] : _GEN_570; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_715 = 8'h8a == _T_10 ? io_in_bits[39:32] : _GEN_571; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_716 = 8'h8b == _T_10 ? io_in_bits[39:32] : _GEN_572; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_717 = 8'h8c == _T_10 ? io_in_bits[39:32] : _GEN_573; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_718 = 8'h8d == _T_10 ? io_in_bits[39:32] : _GEN_574; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_719 = 8'h8e == _T_10 ? io_in_bits[39:32] : _GEN_575; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_720 = 8'h8f == _T_10 ? io_in_bits[39:32] : _GEN_576; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_12 = enqPtr + 8'h5; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_721 = 8'h0 == _T_12 ? io_in_bits[47:40] : _GEN_577; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_722 = 8'h1 == _T_12 ? io_in_bits[47:40] : _GEN_578; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_723 = 8'h2 == _T_12 ? io_in_bits[47:40] : _GEN_579; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_724 = 8'h3 == _T_12 ? io_in_bits[47:40] : _GEN_580; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_725 = 8'h4 == _T_12 ? io_in_bits[47:40] : _GEN_581; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_726 = 8'h5 == _T_12 ? io_in_bits[47:40] : _GEN_582; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_727 = 8'h6 == _T_12 ? io_in_bits[47:40] : _GEN_583; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_728 = 8'h7 == _T_12 ? io_in_bits[47:40] : _GEN_584; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_729 = 8'h8 == _T_12 ? io_in_bits[47:40] : _GEN_585; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_730 = 8'h9 == _T_12 ? io_in_bits[47:40] : _GEN_586; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_731 = 8'ha == _T_12 ? io_in_bits[47:40] : _GEN_587; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_732 = 8'hb == _T_12 ? io_in_bits[47:40] : _GEN_588; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_733 = 8'hc == _T_12 ? io_in_bits[47:40] : _GEN_589; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_734 = 8'hd == _T_12 ? io_in_bits[47:40] : _GEN_590; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_735 = 8'he == _T_12 ? io_in_bits[47:40] : _GEN_591; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_736 = 8'hf == _T_12 ? io_in_bits[47:40] : _GEN_592; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_737 = 8'h10 == _T_12 ? io_in_bits[47:40] : _GEN_593; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_738 = 8'h11 == _T_12 ? io_in_bits[47:40] : _GEN_594; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_739 = 8'h12 == _T_12 ? io_in_bits[47:40] : _GEN_595; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_740 = 8'h13 == _T_12 ? io_in_bits[47:40] : _GEN_596; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_741 = 8'h14 == _T_12 ? io_in_bits[47:40] : _GEN_597; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_742 = 8'h15 == _T_12 ? io_in_bits[47:40] : _GEN_598; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_743 = 8'h16 == _T_12 ? io_in_bits[47:40] : _GEN_599; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_744 = 8'h17 == _T_12 ? io_in_bits[47:40] : _GEN_600; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_745 = 8'h18 == _T_12 ? io_in_bits[47:40] : _GEN_601; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_746 = 8'h19 == _T_12 ? io_in_bits[47:40] : _GEN_602; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_747 = 8'h1a == _T_12 ? io_in_bits[47:40] : _GEN_603; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_748 = 8'h1b == _T_12 ? io_in_bits[47:40] : _GEN_604; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_749 = 8'h1c == _T_12 ? io_in_bits[47:40] : _GEN_605; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_750 = 8'h1d == _T_12 ? io_in_bits[47:40] : _GEN_606; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_751 = 8'h1e == _T_12 ? io_in_bits[47:40] : _GEN_607; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_752 = 8'h1f == _T_12 ? io_in_bits[47:40] : _GEN_608; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_753 = 8'h20 == _T_12 ? io_in_bits[47:40] : _GEN_609; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_754 = 8'h21 == _T_12 ? io_in_bits[47:40] : _GEN_610; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_755 = 8'h22 == _T_12 ? io_in_bits[47:40] : _GEN_611; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_756 = 8'h23 == _T_12 ? io_in_bits[47:40] : _GEN_612; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_757 = 8'h24 == _T_12 ? io_in_bits[47:40] : _GEN_613; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_758 = 8'h25 == _T_12 ? io_in_bits[47:40] : _GEN_614; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_759 = 8'h26 == _T_12 ? io_in_bits[47:40] : _GEN_615; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_760 = 8'h27 == _T_12 ? io_in_bits[47:40] : _GEN_616; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_761 = 8'h28 == _T_12 ? io_in_bits[47:40] : _GEN_617; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_762 = 8'h29 == _T_12 ? io_in_bits[47:40] : _GEN_618; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_763 = 8'h2a == _T_12 ? io_in_bits[47:40] : _GEN_619; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_764 = 8'h2b == _T_12 ? io_in_bits[47:40] : _GEN_620; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_765 = 8'h2c == _T_12 ? io_in_bits[47:40] : _GEN_621; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_766 = 8'h2d == _T_12 ? io_in_bits[47:40] : _GEN_622; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_767 = 8'h2e == _T_12 ? io_in_bits[47:40] : _GEN_623; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_768 = 8'h2f == _T_12 ? io_in_bits[47:40] : _GEN_624; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_769 = 8'h30 == _T_12 ? io_in_bits[47:40] : _GEN_625; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_770 = 8'h31 == _T_12 ? io_in_bits[47:40] : _GEN_626; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_771 = 8'h32 == _T_12 ? io_in_bits[47:40] : _GEN_627; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_772 = 8'h33 == _T_12 ? io_in_bits[47:40] : _GEN_628; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_773 = 8'h34 == _T_12 ? io_in_bits[47:40] : _GEN_629; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_774 = 8'h35 == _T_12 ? io_in_bits[47:40] : _GEN_630; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_775 = 8'h36 == _T_12 ? io_in_bits[47:40] : _GEN_631; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_776 = 8'h37 == _T_12 ? io_in_bits[47:40] : _GEN_632; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_777 = 8'h38 == _T_12 ? io_in_bits[47:40] : _GEN_633; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_778 = 8'h39 == _T_12 ? io_in_bits[47:40] : _GEN_634; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_779 = 8'h3a == _T_12 ? io_in_bits[47:40] : _GEN_635; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_780 = 8'h3b == _T_12 ? io_in_bits[47:40] : _GEN_636; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_781 = 8'h3c == _T_12 ? io_in_bits[47:40] : _GEN_637; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_782 = 8'h3d == _T_12 ? io_in_bits[47:40] : _GEN_638; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_783 = 8'h3e == _T_12 ? io_in_bits[47:40] : _GEN_639; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_784 = 8'h3f == _T_12 ? io_in_bits[47:40] : _GEN_640; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_785 = 8'h40 == _T_12 ? io_in_bits[47:40] : _GEN_641; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_786 = 8'h41 == _T_12 ? io_in_bits[47:40] : _GEN_642; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_787 = 8'h42 == _T_12 ? io_in_bits[47:40] : _GEN_643; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_788 = 8'h43 == _T_12 ? io_in_bits[47:40] : _GEN_644; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_789 = 8'h44 == _T_12 ? io_in_bits[47:40] : _GEN_645; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_790 = 8'h45 == _T_12 ? io_in_bits[47:40] : _GEN_646; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_791 = 8'h46 == _T_12 ? io_in_bits[47:40] : _GEN_647; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_792 = 8'h47 == _T_12 ? io_in_bits[47:40] : _GEN_648; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_793 = 8'h48 == _T_12 ? io_in_bits[47:40] : _GEN_649; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_794 = 8'h49 == _T_12 ? io_in_bits[47:40] : _GEN_650; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_795 = 8'h4a == _T_12 ? io_in_bits[47:40] : _GEN_651; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_796 = 8'h4b == _T_12 ? io_in_bits[47:40] : _GEN_652; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_797 = 8'h4c == _T_12 ? io_in_bits[47:40] : _GEN_653; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_798 = 8'h4d == _T_12 ? io_in_bits[47:40] : _GEN_654; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_799 = 8'h4e == _T_12 ? io_in_bits[47:40] : _GEN_655; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_800 = 8'h4f == _T_12 ? io_in_bits[47:40] : _GEN_656; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_801 = 8'h50 == _T_12 ? io_in_bits[47:40] : _GEN_657; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_802 = 8'h51 == _T_12 ? io_in_bits[47:40] : _GEN_658; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_803 = 8'h52 == _T_12 ? io_in_bits[47:40] : _GEN_659; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_804 = 8'h53 == _T_12 ? io_in_bits[47:40] : _GEN_660; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_805 = 8'h54 == _T_12 ? io_in_bits[47:40] : _GEN_661; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_806 = 8'h55 == _T_12 ? io_in_bits[47:40] : _GEN_662; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_807 = 8'h56 == _T_12 ? io_in_bits[47:40] : _GEN_663; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_808 = 8'h57 == _T_12 ? io_in_bits[47:40] : _GEN_664; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_809 = 8'h58 == _T_12 ? io_in_bits[47:40] : _GEN_665; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_810 = 8'h59 == _T_12 ? io_in_bits[47:40] : _GEN_666; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_811 = 8'h5a == _T_12 ? io_in_bits[47:40] : _GEN_667; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_812 = 8'h5b == _T_12 ? io_in_bits[47:40] : _GEN_668; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_813 = 8'h5c == _T_12 ? io_in_bits[47:40] : _GEN_669; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_814 = 8'h5d == _T_12 ? io_in_bits[47:40] : _GEN_670; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_815 = 8'h5e == _T_12 ? io_in_bits[47:40] : _GEN_671; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_816 = 8'h5f == _T_12 ? io_in_bits[47:40] : _GEN_672; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_817 = 8'h60 == _T_12 ? io_in_bits[47:40] : _GEN_673; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_818 = 8'h61 == _T_12 ? io_in_bits[47:40] : _GEN_674; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_819 = 8'h62 == _T_12 ? io_in_bits[47:40] : _GEN_675; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_820 = 8'h63 == _T_12 ? io_in_bits[47:40] : _GEN_676; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_821 = 8'h64 == _T_12 ? io_in_bits[47:40] : _GEN_677; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_822 = 8'h65 == _T_12 ? io_in_bits[47:40] : _GEN_678; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_823 = 8'h66 == _T_12 ? io_in_bits[47:40] : _GEN_679; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_824 = 8'h67 == _T_12 ? io_in_bits[47:40] : _GEN_680; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_825 = 8'h68 == _T_12 ? io_in_bits[47:40] : _GEN_681; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_826 = 8'h69 == _T_12 ? io_in_bits[47:40] : _GEN_682; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_827 = 8'h6a == _T_12 ? io_in_bits[47:40] : _GEN_683; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_828 = 8'h6b == _T_12 ? io_in_bits[47:40] : _GEN_684; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_829 = 8'h6c == _T_12 ? io_in_bits[47:40] : _GEN_685; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_830 = 8'h6d == _T_12 ? io_in_bits[47:40] : _GEN_686; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_831 = 8'h6e == _T_12 ? io_in_bits[47:40] : _GEN_687; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_832 = 8'h6f == _T_12 ? io_in_bits[47:40] : _GEN_688; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_833 = 8'h70 == _T_12 ? io_in_bits[47:40] : _GEN_689; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_834 = 8'h71 == _T_12 ? io_in_bits[47:40] : _GEN_690; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_835 = 8'h72 == _T_12 ? io_in_bits[47:40] : _GEN_691; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_836 = 8'h73 == _T_12 ? io_in_bits[47:40] : _GEN_692; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_837 = 8'h74 == _T_12 ? io_in_bits[47:40] : _GEN_693; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_838 = 8'h75 == _T_12 ? io_in_bits[47:40] : _GEN_694; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_839 = 8'h76 == _T_12 ? io_in_bits[47:40] : _GEN_695; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_840 = 8'h77 == _T_12 ? io_in_bits[47:40] : _GEN_696; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_841 = 8'h78 == _T_12 ? io_in_bits[47:40] : _GEN_697; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_842 = 8'h79 == _T_12 ? io_in_bits[47:40] : _GEN_698; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_843 = 8'h7a == _T_12 ? io_in_bits[47:40] : _GEN_699; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_844 = 8'h7b == _T_12 ? io_in_bits[47:40] : _GEN_700; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_845 = 8'h7c == _T_12 ? io_in_bits[47:40] : _GEN_701; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_846 = 8'h7d == _T_12 ? io_in_bits[47:40] : _GEN_702; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_847 = 8'h7e == _T_12 ? io_in_bits[47:40] : _GEN_703; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_848 = 8'h7f == _T_12 ? io_in_bits[47:40] : _GEN_704; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_849 = 8'h80 == _T_12 ? io_in_bits[47:40] : _GEN_705; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_850 = 8'h81 == _T_12 ? io_in_bits[47:40] : _GEN_706; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_851 = 8'h82 == _T_12 ? io_in_bits[47:40] : _GEN_707; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_852 = 8'h83 == _T_12 ? io_in_bits[47:40] : _GEN_708; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_853 = 8'h84 == _T_12 ? io_in_bits[47:40] : _GEN_709; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_854 = 8'h85 == _T_12 ? io_in_bits[47:40] : _GEN_710; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_855 = 8'h86 == _T_12 ? io_in_bits[47:40] : _GEN_711; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_856 = 8'h87 == _T_12 ? io_in_bits[47:40] : _GEN_712; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_857 = 8'h88 == _T_12 ? io_in_bits[47:40] : _GEN_713; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_858 = 8'h89 == _T_12 ? io_in_bits[47:40] : _GEN_714; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_859 = 8'h8a == _T_12 ? io_in_bits[47:40] : _GEN_715; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_860 = 8'h8b == _T_12 ? io_in_bits[47:40] : _GEN_716; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_861 = 8'h8c == _T_12 ? io_in_bits[47:40] : _GEN_717; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_862 = 8'h8d == _T_12 ? io_in_bits[47:40] : _GEN_718; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_863 = 8'h8e == _T_12 ? io_in_bits[47:40] : _GEN_719; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_864 = 8'h8f == _T_12 ? io_in_bits[47:40] : _GEN_720; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_14 = enqPtr + 8'h6; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_865 = 8'h0 == _T_14 ? io_in_bits[55:48] : _GEN_721; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_866 = 8'h1 == _T_14 ? io_in_bits[55:48] : _GEN_722; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_867 = 8'h2 == _T_14 ? io_in_bits[55:48] : _GEN_723; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_868 = 8'h3 == _T_14 ? io_in_bits[55:48] : _GEN_724; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_869 = 8'h4 == _T_14 ? io_in_bits[55:48] : _GEN_725; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_870 = 8'h5 == _T_14 ? io_in_bits[55:48] : _GEN_726; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_871 = 8'h6 == _T_14 ? io_in_bits[55:48] : _GEN_727; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_872 = 8'h7 == _T_14 ? io_in_bits[55:48] : _GEN_728; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_873 = 8'h8 == _T_14 ? io_in_bits[55:48] : _GEN_729; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_874 = 8'h9 == _T_14 ? io_in_bits[55:48] : _GEN_730; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_875 = 8'ha == _T_14 ? io_in_bits[55:48] : _GEN_731; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_876 = 8'hb == _T_14 ? io_in_bits[55:48] : _GEN_732; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_877 = 8'hc == _T_14 ? io_in_bits[55:48] : _GEN_733; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_878 = 8'hd == _T_14 ? io_in_bits[55:48] : _GEN_734; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_879 = 8'he == _T_14 ? io_in_bits[55:48] : _GEN_735; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_880 = 8'hf == _T_14 ? io_in_bits[55:48] : _GEN_736; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_881 = 8'h10 == _T_14 ? io_in_bits[55:48] : _GEN_737; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_882 = 8'h11 == _T_14 ? io_in_bits[55:48] : _GEN_738; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_883 = 8'h12 == _T_14 ? io_in_bits[55:48] : _GEN_739; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_884 = 8'h13 == _T_14 ? io_in_bits[55:48] : _GEN_740; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_885 = 8'h14 == _T_14 ? io_in_bits[55:48] : _GEN_741; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_886 = 8'h15 == _T_14 ? io_in_bits[55:48] : _GEN_742; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_887 = 8'h16 == _T_14 ? io_in_bits[55:48] : _GEN_743; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_888 = 8'h17 == _T_14 ? io_in_bits[55:48] : _GEN_744; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_889 = 8'h18 == _T_14 ? io_in_bits[55:48] : _GEN_745; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_890 = 8'h19 == _T_14 ? io_in_bits[55:48] : _GEN_746; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_891 = 8'h1a == _T_14 ? io_in_bits[55:48] : _GEN_747; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_892 = 8'h1b == _T_14 ? io_in_bits[55:48] : _GEN_748; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_893 = 8'h1c == _T_14 ? io_in_bits[55:48] : _GEN_749; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_894 = 8'h1d == _T_14 ? io_in_bits[55:48] : _GEN_750; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_895 = 8'h1e == _T_14 ? io_in_bits[55:48] : _GEN_751; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_896 = 8'h1f == _T_14 ? io_in_bits[55:48] : _GEN_752; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_897 = 8'h20 == _T_14 ? io_in_bits[55:48] : _GEN_753; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_898 = 8'h21 == _T_14 ? io_in_bits[55:48] : _GEN_754; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_899 = 8'h22 == _T_14 ? io_in_bits[55:48] : _GEN_755; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_900 = 8'h23 == _T_14 ? io_in_bits[55:48] : _GEN_756; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_901 = 8'h24 == _T_14 ? io_in_bits[55:48] : _GEN_757; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_902 = 8'h25 == _T_14 ? io_in_bits[55:48] : _GEN_758; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_903 = 8'h26 == _T_14 ? io_in_bits[55:48] : _GEN_759; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_904 = 8'h27 == _T_14 ? io_in_bits[55:48] : _GEN_760; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_905 = 8'h28 == _T_14 ? io_in_bits[55:48] : _GEN_761; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_906 = 8'h29 == _T_14 ? io_in_bits[55:48] : _GEN_762; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_907 = 8'h2a == _T_14 ? io_in_bits[55:48] : _GEN_763; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_908 = 8'h2b == _T_14 ? io_in_bits[55:48] : _GEN_764; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_909 = 8'h2c == _T_14 ? io_in_bits[55:48] : _GEN_765; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_910 = 8'h2d == _T_14 ? io_in_bits[55:48] : _GEN_766; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_911 = 8'h2e == _T_14 ? io_in_bits[55:48] : _GEN_767; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_912 = 8'h2f == _T_14 ? io_in_bits[55:48] : _GEN_768; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_913 = 8'h30 == _T_14 ? io_in_bits[55:48] : _GEN_769; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_914 = 8'h31 == _T_14 ? io_in_bits[55:48] : _GEN_770; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_915 = 8'h32 == _T_14 ? io_in_bits[55:48] : _GEN_771; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_916 = 8'h33 == _T_14 ? io_in_bits[55:48] : _GEN_772; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_917 = 8'h34 == _T_14 ? io_in_bits[55:48] : _GEN_773; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_918 = 8'h35 == _T_14 ? io_in_bits[55:48] : _GEN_774; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_919 = 8'h36 == _T_14 ? io_in_bits[55:48] : _GEN_775; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_920 = 8'h37 == _T_14 ? io_in_bits[55:48] : _GEN_776; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_921 = 8'h38 == _T_14 ? io_in_bits[55:48] : _GEN_777; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_922 = 8'h39 == _T_14 ? io_in_bits[55:48] : _GEN_778; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_923 = 8'h3a == _T_14 ? io_in_bits[55:48] : _GEN_779; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_924 = 8'h3b == _T_14 ? io_in_bits[55:48] : _GEN_780; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_925 = 8'h3c == _T_14 ? io_in_bits[55:48] : _GEN_781; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_926 = 8'h3d == _T_14 ? io_in_bits[55:48] : _GEN_782; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_927 = 8'h3e == _T_14 ? io_in_bits[55:48] : _GEN_783; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_928 = 8'h3f == _T_14 ? io_in_bits[55:48] : _GEN_784; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_929 = 8'h40 == _T_14 ? io_in_bits[55:48] : _GEN_785; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_930 = 8'h41 == _T_14 ? io_in_bits[55:48] : _GEN_786; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_931 = 8'h42 == _T_14 ? io_in_bits[55:48] : _GEN_787; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_932 = 8'h43 == _T_14 ? io_in_bits[55:48] : _GEN_788; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_933 = 8'h44 == _T_14 ? io_in_bits[55:48] : _GEN_789; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_934 = 8'h45 == _T_14 ? io_in_bits[55:48] : _GEN_790; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_935 = 8'h46 == _T_14 ? io_in_bits[55:48] : _GEN_791; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_936 = 8'h47 == _T_14 ? io_in_bits[55:48] : _GEN_792; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_937 = 8'h48 == _T_14 ? io_in_bits[55:48] : _GEN_793; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_938 = 8'h49 == _T_14 ? io_in_bits[55:48] : _GEN_794; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_939 = 8'h4a == _T_14 ? io_in_bits[55:48] : _GEN_795; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_940 = 8'h4b == _T_14 ? io_in_bits[55:48] : _GEN_796; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_941 = 8'h4c == _T_14 ? io_in_bits[55:48] : _GEN_797; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_942 = 8'h4d == _T_14 ? io_in_bits[55:48] : _GEN_798; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_943 = 8'h4e == _T_14 ? io_in_bits[55:48] : _GEN_799; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_944 = 8'h4f == _T_14 ? io_in_bits[55:48] : _GEN_800; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_945 = 8'h50 == _T_14 ? io_in_bits[55:48] : _GEN_801; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_946 = 8'h51 == _T_14 ? io_in_bits[55:48] : _GEN_802; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_947 = 8'h52 == _T_14 ? io_in_bits[55:48] : _GEN_803; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_948 = 8'h53 == _T_14 ? io_in_bits[55:48] : _GEN_804; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_949 = 8'h54 == _T_14 ? io_in_bits[55:48] : _GEN_805; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_950 = 8'h55 == _T_14 ? io_in_bits[55:48] : _GEN_806; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_951 = 8'h56 == _T_14 ? io_in_bits[55:48] : _GEN_807; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_952 = 8'h57 == _T_14 ? io_in_bits[55:48] : _GEN_808; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_953 = 8'h58 == _T_14 ? io_in_bits[55:48] : _GEN_809; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_954 = 8'h59 == _T_14 ? io_in_bits[55:48] : _GEN_810; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_955 = 8'h5a == _T_14 ? io_in_bits[55:48] : _GEN_811; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_956 = 8'h5b == _T_14 ? io_in_bits[55:48] : _GEN_812; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_957 = 8'h5c == _T_14 ? io_in_bits[55:48] : _GEN_813; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_958 = 8'h5d == _T_14 ? io_in_bits[55:48] : _GEN_814; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_959 = 8'h5e == _T_14 ? io_in_bits[55:48] : _GEN_815; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_960 = 8'h5f == _T_14 ? io_in_bits[55:48] : _GEN_816; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_961 = 8'h60 == _T_14 ? io_in_bits[55:48] : _GEN_817; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_962 = 8'h61 == _T_14 ? io_in_bits[55:48] : _GEN_818; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_963 = 8'h62 == _T_14 ? io_in_bits[55:48] : _GEN_819; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_964 = 8'h63 == _T_14 ? io_in_bits[55:48] : _GEN_820; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_965 = 8'h64 == _T_14 ? io_in_bits[55:48] : _GEN_821; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_966 = 8'h65 == _T_14 ? io_in_bits[55:48] : _GEN_822; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_967 = 8'h66 == _T_14 ? io_in_bits[55:48] : _GEN_823; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_968 = 8'h67 == _T_14 ? io_in_bits[55:48] : _GEN_824; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_969 = 8'h68 == _T_14 ? io_in_bits[55:48] : _GEN_825; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_970 = 8'h69 == _T_14 ? io_in_bits[55:48] : _GEN_826; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_971 = 8'h6a == _T_14 ? io_in_bits[55:48] : _GEN_827; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_972 = 8'h6b == _T_14 ? io_in_bits[55:48] : _GEN_828; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_973 = 8'h6c == _T_14 ? io_in_bits[55:48] : _GEN_829; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_974 = 8'h6d == _T_14 ? io_in_bits[55:48] : _GEN_830; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_975 = 8'h6e == _T_14 ? io_in_bits[55:48] : _GEN_831; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_976 = 8'h6f == _T_14 ? io_in_bits[55:48] : _GEN_832; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_977 = 8'h70 == _T_14 ? io_in_bits[55:48] : _GEN_833; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_978 = 8'h71 == _T_14 ? io_in_bits[55:48] : _GEN_834; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_979 = 8'h72 == _T_14 ? io_in_bits[55:48] : _GEN_835; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_980 = 8'h73 == _T_14 ? io_in_bits[55:48] : _GEN_836; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_981 = 8'h74 == _T_14 ? io_in_bits[55:48] : _GEN_837; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_982 = 8'h75 == _T_14 ? io_in_bits[55:48] : _GEN_838; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_983 = 8'h76 == _T_14 ? io_in_bits[55:48] : _GEN_839; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_984 = 8'h77 == _T_14 ? io_in_bits[55:48] : _GEN_840; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_985 = 8'h78 == _T_14 ? io_in_bits[55:48] : _GEN_841; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_986 = 8'h79 == _T_14 ? io_in_bits[55:48] : _GEN_842; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_987 = 8'h7a == _T_14 ? io_in_bits[55:48] : _GEN_843; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_988 = 8'h7b == _T_14 ? io_in_bits[55:48] : _GEN_844; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_989 = 8'h7c == _T_14 ? io_in_bits[55:48] : _GEN_845; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_990 = 8'h7d == _T_14 ? io_in_bits[55:48] : _GEN_846; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_991 = 8'h7e == _T_14 ? io_in_bits[55:48] : _GEN_847; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_992 = 8'h7f == _T_14 ? io_in_bits[55:48] : _GEN_848; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_993 = 8'h80 == _T_14 ? io_in_bits[55:48] : _GEN_849; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_994 = 8'h81 == _T_14 ? io_in_bits[55:48] : _GEN_850; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_995 = 8'h82 == _T_14 ? io_in_bits[55:48] : _GEN_851; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_996 = 8'h83 == _T_14 ? io_in_bits[55:48] : _GEN_852; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_997 = 8'h84 == _T_14 ? io_in_bits[55:48] : _GEN_853; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_998 = 8'h85 == _T_14 ? io_in_bits[55:48] : _GEN_854; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_999 = 8'h86 == _T_14 ? io_in_bits[55:48] : _GEN_855; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1000 = 8'h87 == _T_14 ? io_in_bits[55:48] : _GEN_856; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1001 = 8'h88 == _T_14 ? io_in_bits[55:48] : _GEN_857; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1002 = 8'h89 == _T_14 ? io_in_bits[55:48] : _GEN_858; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1003 = 8'h8a == _T_14 ? io_in_bits[55:48] : _GEN_859; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1004 = 8'h8b == _T_14 ? io_in_bits[55:48] : _GEN_860; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1005 = 8'h8c == _T_14 ? io_in_bits[55:48] : _GEN_861; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1006 = 8'h8d == _T_14 ? io_in_bits[55:48] : _GEN_862; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1007 = 8'h8e == _T_14 ? io_in_bits[55:48] : _GEN_863; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1008 = 8'h8f == _T_14 ? io_in_bits[55:48] : _GEN_864; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_16 = enqPtr + 8'h7; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_1009 = 8'h0 == _T_16 ? io_in_bits[63:56] : _GEN_865; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1010 = 8'h1 == _T_16 ? io_in_bits[63:56] : _GEN_866; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1011 = 8'h2 == _T_16 ? io_in_bits[63:56] : _GEN_867; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1012 = 8'h3 == _T_16 ? io_in_bits[63:56] : _GEN_868; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1013 = 8'h4 == _T_16 ? io_in_bits[63:56] : _GEN_869; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1014 = 8'h5 == _T_16 ? io_in_bits[63:56] : _GEN_870; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1015 = 8'h6 == _T_16 ? io_in_bits[63:56] : _GEN_871; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1016 = 8'h7 == _T_16 ? io_in_bits[63:56] : _GEN_872; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1017 = 8'h8 == _T_16 ? io_in_bits[63:56] : _GEN_873; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1018 = 8'h9 == _T_16 ? io_in_bits[63:56] : _GEN_874; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1019 = 8'ha == _T_16 ? io_in_bits[63:56] : _GEN_875; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1020 = 8'hb == _T_16 ? io_in_bits[63:56] : _GEN_876; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1021 = 8'hc == _T_16 ? io_in_bits[63:56] : _GEN_877; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1022 = 8'hd == _T_16 ? io_in_bits[63:56] : _GEN_878; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1023 = 8'he == _T_16 ? io_in_bits[63:56] : _GEN_879; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1024 = 8'hf == _T_16 ? io_in_bits[63:56] : _GEN_880; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1025 = 8'h10 == _T_16 ? io_in_bits[63:56] : _GEN_881; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1026 = 8'h11 == _T_16 ? io_in_bits[63:56] : _GEN_882; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1027 = 8'h12 == _T_16 ? io_in_bits[63:56] : _GEN_883; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1028 = 8'h13 == _T_16 ? io_in_bits[63:56] : _GEN_884; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1029 = 8'h14 == _T_16 ? io_in_bits[63:56] : _GEN_885; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1030 = 8'h15 == _T_16 ? io_in_bits[63:56] : _GEN_886; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1031 = 8'h16 == _T_16 ? io_in_bits[63:56] : _GEN_887; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1032 = 8'h17 == _T_16 ? io_in_bits[63:56] : _GEN_888; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1033 = 8'h18 == _T_16 ? io_in_bits[63:56] : _GEN_889; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1034 = 8'h19 == _T_16 ? io_in_bits[63:56] : _GEN_890; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1035 = 8'h1a == _T_16 ? io_in_bits[63:56] : _GEN_891; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1036 = 8'h1b == _T_16 ? io_in_bits[63:56] : _GEN_892; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1037 = 8'h1c == _T_16 ? io_in_bits[63:56] : _GEN_893; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1038 = 8'h1d == _T_16 ? io_in_bits[63:56] : _GEN_894; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1039 = 8'h1e == _T_16 ? io_in_bits[63:56] : _GEN_895; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1040 = 8'h1f == _T_16 ? io_in_bits[63:56] : _GEN_896; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1041 = 8'h20 == _T_16 ? io_in_bits[63:56] : _GEN_897; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1042 = 8'h21 == _T_16 ? io_in_bits[63:56] : _GEN_898; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1043 = 8'h22 == _T_16 ? io_in_bits[63:56] : _GEN_899; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1044 = 8'h23 == _T_16 ? io_in_bits[63:56] : _GEN_900; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1045 = 8'h24 == _T_16 ? io_in_bits[63:56] : _GEN_901; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1046 = 8'h25 == _T_16 ? io_in_bits[63:56] : _GEN_902; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1047 = 8'h26 == _T_16 ? io_in_bits[63:56] : _GEN_903; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1048 = 8'h27 == _T_16 ? io_in_bits[63:56] : _GEN_904; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1049 = 8'h28 == _T_16 ? io_in_bits[63:56] : _GEN_905; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1050 = 8'h29 == _T_16 ? io_in_bits[63:56] : _GEN_906; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1051 = 8'h2a == _T_16 ? io_in_bits[63:56] : _GEN_907; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1052 = 8'h2b == _T_16 ? io_in_bits[63:56] : _GEN_908; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1053 = 8'h2c == _T_16 ? io_in_bits[63:56] : _GEN_909; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1054 = 8'h2d == _T_16 ? io_in_bits[63:56] : _GEN_910; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1055 = 8'h2e == _T_16 ? io_in_bits[63:56] : _GEN_911; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1056 = 8'h2f == _T_16 ? io_in_bits[63:56] : _GEN_912; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1057 = 8'h30 == _T_16 ? io_in_bits[63:56] : _GEN_913; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1058 = 8'h31 == _T_16 ? io_in_bits[63:56] : _GEN_914; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1059 = 8'h32 == _T_16 ? io_in_bits[63:56] : _GEN_915; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1060 = 8'h33 == _T_16 ? io_in_bits[63:56] : _GEN_916; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1061 = 8'h34 == _T_16 ? io_in_bits[63:56] : _GEN_917; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1062 = 8'h35 == _T_16 ? io_in_bits[63:56] : _GEN_918; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1063 = 8'h36 == _T_16 ? io_in_bits[63:56] : _GEN_919; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1064 = 8'h37 == _T_16 ? io_in_bits[63:56] : _GEN_920; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1065 = 8'h38 == _T_16 ? io_in_bits[63:56] : _GEN_921; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1066 = 8'h39 == _T_16 ? io_in_bits[63:56] : _GEN_922; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1067 = 8'h3a == _T_16 ? io_in_bits[63:56] : _GEN_923; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1068 = 8'h3b == _T_16 ? io_in_bits[63:56] : _GEN_924; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1069 = 8'h3c == _T_16 ? io_in_bits[63:56] : _GEN_925; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1070 = 8'h3d == _T_16 ? io_in_bits[63:56] : _GEN_926; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1071 = 8'h3e == _T_16 ? io_in_bits[63:56] : _GEN_927; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1072 = 8'h3f == _T_16 ? io_in_bits[63:56] : _GEN_928; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1073 = 8'h40 == _T_16 ? io_in_bits[63:56] : _GEN_929; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1074 = 8'h41 == _T_16 ? io_in_bits[63:56] : _GEN_930; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1075 = 8'h42 == _T_16 ? io_in_bits[63:56] : _GEN_931; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1076 = 8'h43 == _T_16 ? io_in_bits[63:56] : _GEN_932; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1077 = 8'h44 == _T_16 ? io_in_bits[63:56] : _GEN_933; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1078 = 8'h45 == _T_16 ? io_in_bits[63:56] : _GEN_934; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1079 = 8'h46 == _T_16 ? io_in_bits[63:56] : _GEN_935; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1080 = 8'h47 == _T_16 ? io_in_bits[63:56] : _GEN_936; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1081 = 8'h48 == _T_16 ? io_in_bits[63:56] : _GEN_937; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1082 = 8'h49 == _T_16 ? io_in_bits[63:56] : _GEN_938; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1083 = 8'h4a == _T_16 ? io_in_bits[63:56] : _GEN_939; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1084 = 8'h4b == _T_16 ? io_in_bits[63:56] : _GEN_940; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1085 = 8'h4c == _T_16 ? io_in_bits[63:56] : _GEN_941; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1086 = 8'h4d == _T_16 ? io_in_bits[63:56] : _GEN_942; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1087 = 8'h4e == _T_16 ? io_in_bits[63:56] : _GEN_943; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1088 = 8'h4f == _T_16 ? io_in_bits[63:56] : _GEN_944; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1089 = 8'h50 == _T_16 ? io_in_bits[63:56] : _GEN_945; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1090 = 8'h51 == _T_16 ? io_in_bits[63:56] : _GEN_946; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1091 = 8'h52 == _T_16 ? io_in_bits[63:56] : _GEN_947; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1092 = 8'h53 == _T_16 ? io_in_bits[63:56] : _GEN_948; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1093 = 8'h54 == _T_16 ? io_in_bits[63:56] : _GEN_949; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1094 = 8'h55 == _T_16 ? io_in_bits[63:56] : _GEN_950; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1095 = 8'h56 == _T_16 ? io_in_bits[63:56] : _GEN_951; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1096 = 8'h57 == _T_16 ? io_in_bits[63:56] : _GEN_952; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1097 = 8'h58 == _T_16 ? io_in_bits[63:56] : _GEN_953; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1098 = 8'h59 == _T_16 ? io_in_bits[63:56] : _GEN_954; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1099 = 8'h5a == _T_16 ? io_in_bits[63:56] : _GEN_955; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1100 = 8'h5b == _T_16 ? io_in_bits[63:56] : _GEN_956; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1101 = 8'h5c == _T_16 ? io_in_bits[63:56] : _GEN_957; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1102 = 8'h5d == _T_16 ? io_in_bits[63:56] : _GEN_958; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1103 = 8'h5e == _T_16 ? io_in_bits[63:56] : _GEN_959; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1104 = 8'h5f == _T_16 ? io_in_bits[63:56] : _GEN_960; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1105 = 8'h60 == _T_16 ? io_in_bits[63:56] : _GEN_961; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1106 = 8'h61 == _T_16 ? io_in_bits[63:56] : _GEN_962; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1107 = 8'h62 == _T_16 ? io_in_bits[63:56] : _GEN_963; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1108 = 8'h63 == _T_16 ? io_in_bits[63:56] : _GEN_964; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1109 = 8'h64 == _T_16 ? io_in_bits[63:56] : _GEN_965; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1110 = 8'h65 == _T_16 ? io_in_bits[63:56] : _GEN_966; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1111 = 8'h66 == _T_16 ? io_in_bits[63:56] : _GEN_967; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1112 = 8'h67 == _T_16 ? io_in_bits[63:56] : _GEN_968; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1113 = 8'h68 == _T_16 ? io_in_bits[63:56] : _GEN_969; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1114 = 8'h69 == _T_16 ? io_in_bits[63:56] : _GEN_970; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1115 = 8'h6a == _T_16 ? io_in_bits[63:56] : _GEN_971; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1116 = 8'h6b == _T_16 ? io_in_bits[63:56] : _GEN_972; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1117 = 8'h6c == _T_16 ? io_in_bits[63:56] : _GEN_973; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1118 = 8'h6d == _T_16 ? io_in_bits[63:56] : _GEN_974; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1119 = 8'h6e == _T_16 ? io_in_bits[63:56] : _GEN_975; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1120 = 8'h6f == _T_16 ? io_in_bits[63:56] : _GEN_976; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1121 = 8'h70 == _T_16 ? io_in_bits[63:56] : _GEN_977; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1122 = 8'h71 == _T_16 ? io_in_bits[63:56] : _GEN_978; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1123 = 8'h72 == _T_16 ? io_in_bits[63:56] : _GEN_979; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1124 = 8'h73 == _T_16 ? io_in_bits[63:56] : _GEN_980; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1125 = 8'h74 == _T_16 ? io_in_bits[63:56] : _GEN_981; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1126 = 8'h75 == _T_16 ? io_in_bits[63:56] : _GEN_982; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1127 = 8'h76 == _T_16 ? io_in_bits[63:56] : _GEN_983; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1128 = 8'h77 == _T_16 ? io_in_bits[63:56] : _GEN_984; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1129 = 8'h78 == _T_16 ? io_in_bits[63:56] : _GEN_985; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1130 = 8'h79 == _T_16 ? io_in_bits[63:56] : _GEN_986; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1131 = 8'h7a == _T_16 ? io_in_bits[63:56] : _GEN_987; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1132 = 8'h7b == _T_16 ? io_in_bits[63:56] : _GEN_988; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1133 = 8'h7c == _T_16 ? io_in_bits[63:56] : _GEN_989; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1134 = 8'h7d == _T_16 ? io_in_bits[63:56] : _GEN_990; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1135 = 8'h7e == _T_16 ? io_in_bits[63:56] : _GEN_991; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1136 = 8'h7f == _T_16 ? io_in_bits[63:56] : _GEN_992; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1137 = 8'h80 == _T_16 ? io_in_bits[63:56] : _GEN_993; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1138 = 8'h81 == _T_16 ? io_in_bits[63:56] : _GEN_994; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1139 = 8'h82 == _T_16 ? io_in_bits[63:56] : _GEN_995; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1140 = 8'h83 == _T_16 ? io_in_bits[63:56] : _GEN_996; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1141 = 8'h84 == _T_16 ? io_in_bits[63:56] : _GEN_997; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1142 = 8'h85 == _T_16 ? io_in_bits[63:56] : _GEN_998; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1143 = 8'h86 == _T_16 ? io_in_bits[63:56] : _GEN_999; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1144 = 8'h87 == _T_16 ? io_in_bits[63:56] : _GEN_1000; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1145 = 8'h88 == _T_16 ? io_in_bits[63:56] : _GEN_1001; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1146 = 8'h89 == _T_16 ? io_in_bits[63:56] : _GEN_1002; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1147 = 8'h8a == _T_16 ? io_in_bits[63:56] : _GEN_1003; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1148 = 8'h8b == _T_16 ? io_in_bits[63:56] : _GEN_1004; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1149 = 8'h8c == _T_16 ? io_in_bits[63:56] : _GEN_1005; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1150 = 8'h8d == _T_16 ? io_in_bits[63:56] : _GEN_1006; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1151 = 8'h8e == _T_16 ? io_in_bits[63:56] : _GEN_1007; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1152 = 8'h8f == _T_16 ? io_in_bits[63:56] : _GEN_1008; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_18 = enqPtr + 8'h8; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_1153 = 8'h0 == _T_18 ? io_in_bits[71:64] : _GEN_1009; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1154 = 8'h1 == _T_18 ? io_in_bits[71:64] : _GEN_1010; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1155 = 8'h2 == _T_18 ? io_in_bits[71:64] : _GEN_1011; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1156 = 8'h3 == _T_18 ? io_in_bits[71:64] : _GEN_1012; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1157 = 8'h4 == _T_18 ? io_in_bits[71:64] : _GEN_1013; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1158 = 8'h5 == _T_18 ? io_in_bits[71:64] : _GEN_1014; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1159 = 8'h6 == _T_18 ? io_in_bits[71:64] : _GEN_1015; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1160 = 8'h7 == _T_18 ? io_in_bits[71:64] : _GEN_1016; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1161 = 8'h8 == _T_18 ? io_in_bits[71:64] : _GEN_1017; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1162 = 8'h9 == _T_18 ? io_in_bits[71:64] : _GEN_1018; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1163 = 8'ha == _T_18 ? io_in_bits[71:64] : _GEN_1019; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1164 = 8'hb == _T_18 ? io_in_bits[71:64] : _GEN_1020; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1165 = 8'hc == _T_18 ? io_in_bits[71:64] : _GEN_1021; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1166 = 8'hd == _T_18 ? io_in_bits[71:64] : _GEN_1022; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1167 = 8'he == _T_18 ? io_in_bits[71:64] : _GEN_1023; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1168 = 8'hf == _T_18 ? io_in_bits[71:64] : _GEN_1024; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1169 = 8'h10 == _T_18 ? io_in_bits[71:64] : _GEN_1025; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1170 = 8'h11 == _T_18 ? io_in_bits[71:64] : _GEN_1026; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1171 = 8'h12 == _T_18 ? io_in_bits[71:64] : _GEN_1027; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1172 = 8'h13 == _T_18 ? io_in_bits[71:64] : _GEN_1028; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1173 = 8'h14 == _T_18 ? io_in_bits[71:64] : _GEN_1029; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1174 = 8'h15 == _T_18 ? io_in_bits[71:64] : _GEN_1030; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1175 = 8'h16 == _T_18 ? io_in_bits[71:64] : _GEN_1031; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1176 = 8'h17 == _T_18 ? io_in_bits[71:64] : _GEN_1032; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1177 = 8'h18 == _T_18 ? io_in_bits[71:64] : _GEN_1033; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1178 = 8'h19 == _T_18 ? io_in_bits[71:64] : _GEN_1034; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1179 = 8'h1a == _T_18 ? io_in_bits[71:64] : _GEN_1035; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1180 = 8'h1b == _T_18 ? io_in_bits[71:64] : _GEN_1036; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1181 = 8'h1c == _T_18 ? io_in_bits[71:64] : _GEN_1037; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1182 = 8'h1d == _T_18 ? io_in_bits[71:64] : _GEN_1038; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1183 = 8'h1e == _T_18 ? io_in_bits[71:64] : _GEN_1039; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1184 = 8'h1f == _T_18 ? io_in_bits[71:64] : _GEN_1040; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1185 = 8'h20 == _T_18 ? io_in_bits[71:64] : _GEN_1041; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1186 = 8'h21 == _T_18 ? io_in_bits[71:64] : _GEN_1042; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1187 = 8'h22 == _T_18 ? io_in_bits[71:64] : _GEN_1043; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1188 = 8'h23 == _T_18 ? io_in_bits[71:64] : _GEN_1044; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1189 = 8'h24 == _T_18 ? io_in_bits[71:64] : _GEN_1045; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1190 = 8'h25 == _T_18 ? io_in_bits[71:64] : _GEN_1046; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1191 = 8'h26 == _T_18 ? io_in_bits[71:64] : _GEN_1047; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1192 = 8'h27 == _T_18 ? io_in_bits[71:64] : _GEN_1048; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1193 = 8'h28 == _T_18 ? io_in_bits[71:64] : _GEN_1049; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1194 = 8'h29 == _T_18 ? io_in_bits[71:64] : _GEN_1050; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1195 = 8'h2a == _T_18 ? io_in_bits[71:64] : _GEN_1051; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1196 = 8'h2b == _T_18 ? io_in_bits[71:64] : _GEN_1052; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1197 = 8'h2c == _T_18 ? io_in_bits[71:64] : _GEN_1053; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1198 = 8'h2d == _T_18 ? io_in_bits[71:64] : _GEN_1054; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1199 = 8'h2e == _T_18 ? io_in_bits[71:64] : _GEN_1055; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1200 = 8'h2f == _T_18 ? io_in_bits[71:64] : _GEN_1056; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1201 = 8'h30 == _T_18 ? io_in_bits[71:64] : _GEN_1057; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1202 = 8'h31 == _T_18 ? io_in_bits[71:64] : _GEN_1058; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1203 = 8'h32 == _T_18 ? io_in_bits[71:64] : _GEN_1059; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1204 = 8'h33 == _T_18 ? io_in_bits[71:64] : _GEN_1060; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1205 = 8'h34 == _T_18 ? io_in_bits[71:64] : _GEN_1061; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1206 = 8'h35 == _T_18 ? io_in_bits[71:64] : _GEN_1062; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1207 = 8'h36 == _T_18 ? io_in_bits[71:64] : _GEN_1063; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1208 = 8'h37 == _T_18 ? io_in_bits[71:64] : _GEN_1064; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1209 = 8'h38 == _T_18 ? io_in_bits[71:64] : _GEN_1065; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1210 = 8'h39 == _T_18 ? io_in_bits[71:64] : _GEN_1066; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1211 = 8'h3a == _T_18 ? io_in_bits[71:64] : _GEN_1067; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1212 = 8'h3b == _T_18 ? io_in_bits[71:64] : _GEN_1068; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1213 = 8'h3c == _T_18 ? io_in_bits[71:64] : _GEN_1069; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1214 = 8'h3d == _T_18 ? io_in_bits[71:64] : _GEN_1070; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1215 = 8'h3e == _T_18 ? io_in_bits[71:64] : _GEN_1071; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1216 = 8'h3f == _T_18 ? io_in_bits[71:64] : _GEN_1072; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1217 = 8'h40 == _T_18 ? io_in_bits[71:64] : _GEN_1073; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1218 = 8'h41 == _T_18 ? io_in_bits[71:64] : _GEN_1074; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1219 = 8'h42 == _T_18 ? io_in_bits[71:64] : _GEN_1075; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1220 = 8'h43 == _T_18 ? io_in_bits[71:64] : _GEN_1076; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1221 = 8'h44 == _T_18 ? io_in_bits[71:64] : _GEN_1077; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1222 = 8'h45 == _T_18 ? io_in_bits[71:64] : _GEN_1078; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1223 = 8'h46 == _T_18 ? io_in_bits[71:64] : _GEN_1079; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1224 = 8'h47 == _T_18 ? io_in_bits[71:64] : _GEN_1080; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1225 = 8'h48 == _T_18 ? io_in_bits[71:64] : _GEN_1081; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1226 = 8'h49 == _T_18 ? io_in_bits[71:64] : _GEN_1082; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1227 = 8'h4a == _T_18 ? io_in_bits[71:64] : _GEN_1083; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1228 = 8'h4b == _T_18 ? io_in_bits[71:64] : _GEN_1084; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1229 = 8'h4c == _T_18 ? io_in_bits[71:64] : _GEN_1085; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1230 = 8'h4d == _T_18 ? io_in_bits[71:64] : _GEN_1086; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1231 = 8'h4e == _T_18 ? io_in_bits[71:64] : _GEN_1087; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1232 = 8'h4f == _T_18 ? io_in_bits[71:64] : _GEN_1088; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1233 = 8'h50 == _T_18 ? io_in_bits[71:64] : _GEN_1089; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1234 = 8'h51 == _T_18 ? io_in_bits[71:64] : _GEN_1090; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1235 = 8'h52 == _T_18 ? io_in_bits[71:64] : _GEN_1091; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1236 = 8'h53 == _T_18 ? io_in_bits[71:64] : _GEN_1092; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1237 = 8'h54 == _T_18 ? io_in_bits[71:64] : _GEN_1093; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1238 = 8'h55 == _T_18 ? io_in_bits[71:64] : _GEN_1094; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1239 = 8'h56 == _T_18 ? io_in_bits[71:64] : _GEN_1095; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1240 = 8'h57 == _T_18 ? io_in_bits[71:64] : _GEN_1096; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1241 = 8'h58 == _T_18 ? io_in_bits[71:64] : _GEN_1097; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1242 = 8'h59 == _T_18 ? io_in_bits[71:64] : _GEN_1098; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1243 = 8'h5a == _T_18 ? io_in_bits[71:64] : _GEN_1099; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1244 = 8'h5b == _T_18 ? io_in_bits[71:64] : _GEN_1100; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1245 = 8'h5c == _T_18 ? io_in_bits[71:64] : _GEN_1101; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1246 = 8'h5d == _T_18 ? io_in_bits[71:64] : _GEN_1102; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1247 = 8'h5e == _T_18 ? io_in_bits[71:64] : _GEN_1103; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1248 = 8'h5f == _T_18 ? io_in_bits[71:64] : _GEN_1104; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1249 = 8'h60 == _T_18 ? io_in_bits[71:64] : _GEN_1105; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1250 = 8'h61 == _T_18 ? io_in_bits[71:64] : _GEN_1106; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1251 = 8'h62 == _T_18 ? io_in_bits[71:64] : _GEN_1107; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1252 = 8'h63 == _T_18 ? io_in_bits[71:64] : _GEN_1108; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1253 = 8'h64 == _T_18 ? io_in_bits[71:64] : _GEN_1109; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1254 = 8'h65 == _T_18 ? io_in_bits[71:64] : _GEN_1110; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1255 = 8'h66 == _T_18 ? io_in_bits[71:64] : _GEN_1111; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1256 = 8'h67 == _T_18 ? io_in_bits[71:64] : _GEN_1112; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1257 = 8'h68 == _T_18 ? io_in_bits[71:64] : _GEN_1113; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1258 = 8'h69 == _T_18 ? io_in_bits[71:64] : _GEN_1114; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1259 = 8'h6a == _T_18 ? io_in_bits[71:64] : _GEN_1115; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1260 = 8'h6b == _T_18 ? io_in_bits[71:64] : _GEN_1116; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1261 = 8'h6c == _T_18 ? io_in_bits[71:64] : _GEN_1117; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1262 = 8'h6d == _T_18 ? io_in_bits[71:64] : _GEN_1118; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1263 = 8'h6e == _T_18 ? io_in_bits[71:64] : _GEN_1119; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1264 = 8'h6f == _T_18 ? io_in_bits[71:64] : _GEN_1120; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1265 = 8'h70 == _T_18 ? io_in_bits[71:64] : _GEN_1121; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1266 = 8'h71 == _T_18 ? io_in_bits[71:64] : _GEN_1122; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1267 = 8'h72 == _T_18 ? io_in_bits[71:64] : _GEN_1123; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1268 = 8'h73 == _T_18 ? io_in_bits[71:64] : _GEN_1124; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1269 = 8'h74 == _T_18 ? io_in_bits[71:64] : _GEN_1125; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1270 = 8'h75 == _T_18 ? io_in_bits[71:64] : _GEN_1126; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1271 = 8'h76 == _T_18 ? io_in_bits[71:64] : _GEN_1127; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1272 = 8'h77 == _T_18 ? io_in_bits[71:64] : _GEN_1128; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1273 = 8'h78 == _T_18 ? io_in_bits[71:64] : _GEN_1129; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1274 = 8'h79 == _T_18 ? io_in_bits[71:64] : _GEN_1130; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1275 = 8'h7a == _T_18 ? io_in_bits[71:64] : _GEN_1131; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1276 = 8'h7b == _T_18 ? io_in_bits[71:64] : _GEN_1132; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1277 = 8'h7c == _T_18 ? io_in_bits[71:64] : _GEN_1133; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1278 = 8'h7d == _T_18 ? io_in_bits[71:64] : _GEN_1134; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1279 = 8'h7e == _T_18 ? io_in_bits[71:64] : _GEN_1135; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1280 = 8'h7f == _T_18 ? io_in_bits[71:64] : _GEN_1136; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1281 = 8'h80 == _T_18 ? io_in_bits[71:64] : _GEN_1137; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1282 = 8'h81 == _T_18 ? io_in_bits[71:64] : _GEN_1138; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1283 = 8'h82 == _T_18 ? io_in_bits[71:64] : _GEN_1139; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1284 = 8'h83 == _T_18 ? io_in_bits[71:64] : _GEN_1140; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1285 = 8'h84 == _T_18 ? io_in_bits[71:64] : _GEN_1141; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1286 = 8'h85 == _T_18 ? io_in_bits[71:64] : _GEN_1142; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1287 = 8'h86 == _T_18 ? io_in_bits[71:64] : _GEN_1143; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1288 = 8'h87 == _T_18 ? io_in_bits[71:64] : _GEN_1144; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1289 = 8'h88 == _T_18 ? io_in_bits[71:64] : _GEN_1145; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1290 = 8'h89 == _T_18 ? io_in_bits[71:64] : _GEN_1146; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1291 = 8'h8a == _T_18 ? io_in_bits[71:64] : _GEN_1147; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1292 = 8'h8b == _T_18 ? io_in_bits[71:64] : _GEN_1148; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1293 = 8'h8c == _T_18 ? io_in_bits[71:64] : _GEN_1149; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1294 = 8'h8d == _T_18 ? io_in_bits[71:64] : _GEN_1150; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1295 = 8'h8e == _T_18 ? io_in_bits[71:64] : _GEN_1151; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1296 = 8'h8f == _T_18 ? io_in_bits[71:64] : _GEN_1152; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_20 = enqPtr + 8'h9; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_1297 = 8'h0 == _T_20 ? io_in_bits[79:72] : _GEN_1153; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1298 = 8'h1 == _T_20 ? io_in_bits[79:72] : _GEN_1154; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1299 = 8'h2 == _T_20 ? io_in_bits[79:72] : _GEN_1155; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1300 = 8'h3 == _T_20 ? io_in_bits[79:72] : _GEN_1156; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1301 = 8'h4 == _T_20 ? io_in_bits[79:72] : _GEN_1157; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1302 = 8'h5 == _T_20 ? io_in_bits[79:72] : _GEN_1158; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1303 = 8'h6 == _T_20 ? io_in_bits[79:72] : _GEN_1159; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1304 = 8'h7 == _T_20 ? io_in_bits[79:72] : _GEN_1160; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1305 = 8'h8 == _T_20 ? io_in_bits[79:72] : _GEN_1161; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1306 = 8'h9 == _T_20 ? io_in_bits[79:72] : _GEN_1162; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1307 = 8'ha == _T_20 ? io_in_bits[79:72] : _GEN_1163; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1308 = 8'hb == _T_20 ? io_in_bits[79:72] : _GEN_1164; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1309 = 8'hc == _T_20 ? io_in_bits[79:72] : _GEN_1165; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1310 = 8'hd == _T_20 ? io_in_bits[79:72] : _GEN_1166; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1311 = 8'he == _T_20 ? io_in_bits[79:72] : _GEN_1167; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1312 = 8'hf == _T_20 ? io_in_bits[79:72] : _GEN_1168; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1313 = 8'h10 == _T_20 ? io_in_bits[79:72] : _GEN_1169; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1314 = 8'h11 == _T_20 ? io_in_bits[79:72] : _GEN_1170; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1315 = 8'h12 == _T_20 ? io_in_bits[79:72] : _GEN_1171; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1316 = 8'h13 == _T_20 ? io_in_bits[79:72] : _GEN_1172; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1317 = 8'h14 == _T_20 ? io_in_bits[79:72] : _GEN_1173; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1318 = 8'h15 == _T_20 ? io_in_bits[79:72] : _GEN_1174; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1319 = 8'h16 == _T_20 ? io_in_bits[79:72] : _GEN_1175; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1320 = 8'h17 == _T_20 ? io_in_bits[79:72] : _GEN_1176; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1321 = 8'h18 == _T_20 ? io_in_bits[79:72] : _GEN_1177; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1322 = 8'h19 == _T_20 ? io_in_bits[79:72] : _GEN_1178; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1323 = 8'h1a == _T_20 ? io_in_bits[79:72] : _GEN_1179; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1324 = 8'h1b == _T_20 ? io_in_bits[79:72] : _GEN_1180; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1325 = 8'h1c == _T_20 ? io_in_bits[79:72] : _GEN_1181; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1326 = 8'h1d == _T_20 ? io_in_bits[79:72] : _GEN_1182; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1327 = 8'h1e == _T_20 ? io_in_bits[79:72] : _GEN_1183; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1328 = 8'h1f == _T_20 ? io_in_bits[79:72] : _GEN_1184; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1329 = 8'h20 == _T_20 ? io_in_bits[79:72] : _GEN_1185; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1330 = 8'h21 == _T_20 ? io_in_bits[79:72] : _GEN_1186; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1331 = 8'h22 == _T_20 ? io_in_bits[79:72] : _GEN_1187; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1332 = 8'h23 == _T_20 ? io_in_bits[79:72] : _GEN_1188; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1333 = 8'h24 == _T_20 ? io_in_bits[79:72] : _GEN_1189; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1334 = 8'h25 == _T_20 ? io_in_bits[79:72] : _GEN_1190; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1335 = 8'h26 == _T_20 ? io_in_bits[79:72] : _GEN_1191; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1336 = 8'h27 == _T_20 ? io_in_bits[79:72] : _GEN_1192; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1337 = 8'h28 == _T_20 ? io_in_bits[79:72] : _GEN_1193; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1338 = 8'h29 == _T_20 ? io_in_bits[79:72] : _GEN_1194; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1339 = 8'h2a == _T_20 ? io_in_bits[79:72] : _GEN_1195; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1340 = 8'h2b == _T_20 ? io_in_bits[79:72] : _GEN_1196; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1341 = 8'h2c == _T_20 ? io_in_bits[79:72] : _GEN_1197; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1342 = 8'h2d == _T_20 ? io_in_bits[79:72] : _GEN_1198; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1343 = 8'h2e == _T_20 ? io_in_bits[79:72] : _GEN_1199; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1344 = 8'h2f == _T_20 ? io_in_bits[79:72] : _GEN_1200; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1345 = 8'h30 == _T_20 ? io_in_bits[79:72] : _GEN_1201; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1346 = 8'h31 == _T_20 ? io_in_bits[79:72] : _GEN_1202; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1347 = 8'h32 == _T_20 ? io_in_bits[79:72] : _GEN_1203; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1348 = 8'h33 == _T_20 ? io_in_bits[79:72] : _GEN_1204; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1349 = 8'h34 == _T_20 ? io_in_bits[79:72] : _GEN_1205; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1350 = 8'h35 == _T_20 ? io_in_bits[79:72] : _GEN_1206; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1351 = 8'h36 == _T_20 ? io_in_bits[79:72] : _GEN_1207; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1352 = 8'h37 == _T_20 ? io_in_bits[79:72] : _GEN_1208; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1353 = 8'h38 == _T_20 ? io_in_bits[79:72] : _GEN_1209; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1354 = 8'h39 == _T_20 ? io_in_bits[79:72] : _GEN_1210; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1355 = 8'h3a == _T_20 ? io_in_bits[79:72] : _GEN_1211; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1356 = 8'h3b == _T_20 ? io_in_bits[79:72] : _GEN_1212; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1357 = 8'h3c == _T_20 ? io_in_bits[79:72] : _GEN_1213; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1358 = 8'h3d == _T_20 ? io_in_bits[79:72] : _GEN_1214; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1359 = 8'h3e == _T_20 ? io_in_bits[79:72] : _GEN_1215; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1360 = 8'h3f == _T_20 ? io_in_bits[79:72] : _GEN_1216; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1361 = 8'h40 == _T_20 ? io_in_bits[79:72] : _GEN_1217; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1362 = 8'h41 == _T_20 ? io_in_bits[79:72] : _GEN_1218; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1363 = 8'h42 == _T_20 ? io_in_bits[79:72] : _GEN_1219; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1364 = 8'h43 == _T_20 ? io_in_bits[79:72] : _GEN_1220; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1365 = 8'h44 == _T_20 ? io_in_bits[79:72] : _GEN_1221; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1366 = 8'h45 == _T_20 ? io_in_bits[79:72] : _GEN_1222; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1367 = 8'h46 == _T_20 ? io_in_bits[79:72] : _GEN_1223; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1368 = 8'h47 == _T_20 ? io_in_bits[79:72] : _GEN_1224; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1369 = 8'h48 == _T_20 ? io_in_bits[79:72] : _GEN_1225; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1370 = 8'h49 == _T_20 ? io_in_bits[79:72] : _GEN_1226; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1371 = 8'h4a == _T_20 ? io_in_bits[79:72] : _GEN_1227; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1372 = 8'h4b == _T_20 ? io_in_bits[79:72] : _GEN_1228; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1373 = 8'h4c == _T_20 ? io_in_bits[79:72] : _GEN_1229; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1374 = 8'h4d == _T_20 ? io_in_bits[79:72] : _GEN_1230; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1375 = 8'h4e == _T_20 ? io_in_bits[79:72] : _GEN_1231; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1376 = 8'h4f == _T_20 ? io_in_bits[79:72] : _GEN_1232; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1377 = 8'h50 == _T_20 ? io_in_bits[79:72] : _GEN_1233; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1378 = 8'h51 == _T_20 ? io_in_bits[79:72] : _GEN_1234; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1379 = 8'h52 == _T_20 ? io_in_bits[79:72] : _GEN_1235; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1380 = 8'h53 == _T_20 ? io_in_bits[79:72] : _GEN_1236; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1381 = 8'h54 == _T_20 ? io_in_bits[79:72] : _GEN_1237; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1382 = 8'h55 == _T_20 ? io_in_bits[79:72] : _GEN_1238; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1383 = 8'h56 == _T_20 ? io_in_bits[79:72] : _GEN_1239; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1384 = 8'h57 == _T_20 ? io_in_bits[79:72] : _GEN_1240; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1385 = 8'h58 == _T_20 ? io_in_bits[79:72] : _GEN_1241; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1386 = 8'h59 == _T_20 ? io_in_bits[79:72] : _GEN_1242; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1387 = 8'h5a == _T_20 ? io_in_bits[79:72] : _GEN_1243; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1388 = 8'h5b == _T_20 ? io_in_bits[79:72] : _GEN_1244; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1389 = 8'h5c == _T_20 ? io_in_bits[79:72] : _GEN_1245; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1390 = 8'h5d == _T_20 ? io_in_bits[79:72] : _GEN_1246; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1391 = 8'h5e == _T_20 ? io_in_bits[79:72] : _GEN_1247; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1392 = 8'h5f == _T_20 ? io_in_bits[79:72] : _GEN_1248; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1393 = 8'h60 == _T_20 ? io_in_bits[79:72] : _GEN_1249; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1394 = 8'h61 == _T_20 ? io_in_bits[79:72] : _GEN_1250; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1395 = 8'h62 == _T_20 ? io_in_bits[79:72] : _GEN_1251; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1396 = 8'h63 == _T_20 ? io_in_bits[79:72] : _GEN_1252; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1397 = 8'h64 == _T_20 ? io_in_bits[79:72] : _GEN_1253; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1398 = 8'h65 == _T_20 ? io_in_bits[79:72] : _GEN_1254; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1399 = 8'h66 == _T_20 ? io_in_bits[79:72] : _GEN_1255; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1400 = 8'h67 == _T_20 ? io_in_bits[79:72] : _GEN_1256; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1401 = 8'h68 == _T_20 ? io_in_bits[79:72] : _GEN_1257; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1402 = 8'h69 == _T_20 ? io_in_bits[79:72] : _GEN_1258; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1403 = 8'h6a == _T_20 ? io_in_bits[79:72] : _GEN_1259; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1404 = 8'h6b == _T_20 ? io_in_bits[79:72] : _GEN_1260; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1405 = 8'h6c == _T_20 ? io_in_bits[79:72] : _GEN_1261; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1406 = 8'h6d == _T_20 ? io_in_bits[79:72] : _GEN_1262; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1407 = 8'h6e == _T_20 ? io_in_bits[79:72] : _GEN_1263; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1408 = 8'h6f == _T_20 ? io_in_bits[79:72] : _GEN_1264; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1409 = 8'h70 == _T_20 ? io_in_bits[79:72] : _GEN_1265; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1410 = 8'h71 == _T_20 ? io_in_bits[79:72] : _GEN_1266; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1411 = 8'h72 == _T_20 ? io_in_bits[79:72] : _GEN_1267; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1412 = 8'h73 == _T_20 ? io_in_bits[79:72] : _GEN_1268; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1413 = 8'h74 == _T_20 ? io_in_bits[79:72] : _GEN_1269; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1414 = 8'h75 == _T_20 ? io_in_bits[79:72] : _GEN_1270; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1415 = 8'h76 == _T_20 ? io_in_bits[79:72] : _GEN_1271; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1416 = 8'h77 == _T_20 ? io_in_bits[79:72] : _GEN_1272; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1417 = 8'h78 == _T_20 ? io_in_bits[79:72] : _GEN_1273; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1418 = 8'h79 == _T_20 ? io_in_bits[79:72] : _GEN_1274; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1419 = 8'h7a == _T_20 ? io_in_bits[79:72] : _GEN_1275; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1420 = 8'h7b == _T_20 ? io_in_bits[79:72] : _GEN_1276; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1421 = 8'h7c == _T_20 ? io_in_bits[79:72] : _GEN_1277; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1422 = 8'h7d == _T_20 ? io_in_bits[79:72] : _GEN_1278; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1423 = 8'h7e == _T_20 ? io_in_bits[79:72] : _GEN_1279; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1424 = 8'h7f == _T_20 ? io_in_bits[79:72] : _GEN_1280; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1425 = 8'h80 == _T_20 ? io_in_bits[79:72] : _GEN_1281; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1426 = 8'h81 == _T_20 ? io_in_bits[79:72] : _GEN_1282; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1427 = 8'h82 == _T_20 ? io_in_bits[79:72] : _GEN_1283; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1428 = 8'h83 == _T_20 ? io_in_bits[79:72] : _GEN_1284; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1429 = 8'h84 == _T_20 ? io_in_bits[79:72] : _GEN_1285; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1430 = 8'h85 == _T_20 ? io_in_bits[79:72] : _GEN_1286; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1431 = 8'h86 == _T_20 ? io_in_bits[79:72] : _GEN_1287; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1432 = 8'h87 == _T_20 ? io_in_bits[79:72] : _GEN_1288; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1433 = 8'h88 == _T_20 ? io_in_bits[79:72] : _GEN_1289; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1434 = 8'h89 == _T_20 ? io_in_bits[79:72] : _GEN_1290; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1435 = 8'h8a == _T_20 ? io_in_bits[79:72] : _GEN_1291; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1436 = 8'h8b == _T_20 ? io_in_bits[79:72] : _GEN_1292; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1437 = 8'h8c == _T_20 ? io_in_bits[79:72] : _GEN_1293; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1438 = 8'h8d == _T_20 ? io_in_bits[79:72] : _GEN_1294; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1439 = 8'h8e == _T_20 ? io_in_bits[79:72] : _GEN_1295; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1440 = 8'h8f == _T_20 ? io_in_bits[79:72] : _GEN_1296; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_22 = enqPtr + 8'ha; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_1441 = 8'h0 == _T_22 ? io_in_bits[87:80] : _GEN_1297; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1442 = 8'h1 == _T_22 ? io_in_bits[87:80] : _GEN_1298; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1443 = 8'h2 == _T_22 ? io_in_bits[87:80] : _GEN_1299; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1444 = 8'h3 == _T_22 ? io_in_bits[87:80] : _GEN_1300; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1445 = 8'h4 == _T_22 ? io_in_bits[87:80] : _GEN_1301; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1446 = 8'h5 == _T_22 ? io_in_bits[87:80] : _GEN_1302; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1447 = 8'h6 == _T_22 ? io_in_bits[87:80] : _GEN_1303; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1448 = 8'h7 == _T_22 ? io_in_bits[87:80] : _GEN_1304; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1449 = 8'h8 == _T_22 ? io_in_bits[87:80] : _GEN_1305; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1450 = 8'h9 == _T_22 ? io_in_bits[87:80] : _GEN_1306; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1451 = 8'ha == _T_22 ? io_in_bits[87:80] : _GEN_1307; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1452 = 8'hb == _T_22 ? io_in_bits[87:80] : _GEN_1308; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1453 = 8'hc == _T_22 ? io_in_bits[87:80] : _GEN_1309; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1454 = 8'hd == _T_22 ? io_in_bits[87:80] : _GEN_1310; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1455 = 8'he == _T_22 ? io_in_bits[87:80] : _GEN_1311; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1456 = 8'hf == _T_22 ? io_in_bits[87:80] : _GEN_1312; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1457 = 8'h10 == _T_22 ? io_in_bits[87:80] : _GEN_1313; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1458 = 8'h11 == _T_22 ? io_in_bits[87:80] : _GEN_1314; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1459 = 8'h12 == _T_22 ? io_in_bits[87:80] : _GEN_1315; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1460 = 8'h13 == _T_22 ? io_in_bits[87:80] : _GEN_1316; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1461 = 8'h14 == _T_22 ? io_in_bits[87:80] : _GEN_1317; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1462 = 8'h15 == _T_22 ? io_in_bits[87:80] : _GEN_1318; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1463 = 8'h16 == _T_22 ? io_in_bits[87:80] : _GEN_1319; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1464 = 8'h17 == _T_22 ? io_in_bits[87:80] : _GEN_1320; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1465 = 8'h18 == _T_22 ? io_in_bits[87:80] : _GEN_1321; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1466 = 8'h19 == _T_22 ? io_in_bits[87:80] : _GEN_1322; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1467 = 8'h1a == _T_22 ? io_in_bits[87:80] : _GEN_1323; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1468 = 8'h1b == _T_22 ? io_in_bits[87:80] : _GEN_1324; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1469 = 8'h1c == _T_22 ? io_in_bits[87:80] : _GEN_1325; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1470 = 8'h1d == _T_22 ? io_in_bits[87:80] : _GEN_1326; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1471 = 8'h1e == _T_22 ? io_in_bits[87:80] : _GEN_1327; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1472 = 8'h1f == _T_22 ? io_in_bits[87:80] : _GEN_1328; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1473 = 8'h20 == _T_22 ? io_in_bits[87:80] : _GEN_1329; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1474 = 8'h21 == _T_22 ? io_in_bits[87:80] : _GEN_1330; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1475 = 8'h22 == _T_22 ? io_in_bits[87:80] : _GEN_1331; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1476 = 8'h23 == _T_22 ? io_in_bits[87:80] : _GEN_1332; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1477 = 8'h24 == _T_22 ? io_in_bits[87:80] : _GEN_1333; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1478 = 8'h25 == _T_22 ? io_in_bits[87:80] : _GEN_1334; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1479 = 8'h26 == _T_22 ? io_in_bits[87:80] : _GEN_1335; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1480 = 8'h27 == _T_22 ? io_in_bits[87:80] : _GEN_1336; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1481 = 8'h28 == _T_22 ? io_in_bits[87:80] : _GEN_1337; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1482 = 8'h29 == _T_22 ? io_in_bits[87:80] : _GEN_1338; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1483 = 8'h2a == _T_22 ? io_in_bits[87:80] : _GEN_1339; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1484 = 8'h2b == _T_22 ? io_in_bits[87:80] : _GEN_1340; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1485 = 8'h2c == _T_22 ? io_in_bits[87:80] : _GEN_1341; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1486 = 8'h2d == _T_22 ? io_in_bits[87:80] : _GEN_1342; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1487 = 8'h2e == _T_22 ? io_in_bits[87:80] : _GEN_1343; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1488 = 8'h2f == _T_22 ? io_in_bits[87:80] : _GEN_1344; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1489 = 8'h30 == _T_22 ? io_in_bits[87:80] : _GEN_1345; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1490 = 8'h31 == _T_22 ? io_in_bits[87:80] : _GEN_1346; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1491 = 8'h32 == _T_22 ? io_in_bits[87:80] : _GEN_1347; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1492 = 8'h33 == _T_22 ? io_in_bits[87:80] : _GEN_1348; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1493 = 8'h34 == _T_22 ? io_in_bits[87:80] : _GEN_1349; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1494 = 8'h35 == _T_22 ? io_in_bits[87:80] : _GEN_1350; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1495 = 8'h36 == _T_22 ? io_in_bits[87:80] : _GEN_1351; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1496 = 8'h37 == _T_22 ? io_in_bits[87:80] : _GEN_1352; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1497 = 8'h38 == _T_22 ? io_in_bits[87:80] : _GEN_1353; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1498 = 8'h39 == _T_22 ? io_in_bits[87:80] : _GEN_1354; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1499 = 8'h3a == _T_22 ? io_in_bits[87:80] : _GEN_1355; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1500 = 8'h3b == _T_22 ? io_in_bits[87:80] : _GEN_1356; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1501 = 8'h3c == _T_22 ? io_in_bits[87:80] : _GEN_1357; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1502 = 8'h3d == _T_22 ? io_in_bits[87:80] : _GEN_1358; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1503 = 8'h3e == _T_22 ? io_in_bits[87:80] : _GEN_1359; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1504 = 8'h3f == _T_22 ? io_in_bits[87:80] : _GEN_1360; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1505 = 8'h40 == _T_22 ? io_in_bits[87:80] : _GEN_1361; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1506 = 8'h41 == _T_22 ? io_in_bits[87:80] : _GEN_1362; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1507 = 8'h42 == _T_22 ? io_in_bits[87:80] : _GEN_1363; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1508 = 8'h43 == _T_22 ? io_in_bits[87:80] : _GEN_1364; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1509 = 8'h44 == _T_22 ? io_in_bits[87:80] : _GEN_1365; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1510 = 8'h45 == _T_22 ? io_in_bits[87:80] : _GEN_1366; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1511 = 8'h46 == _T_22 ? io_in_bits[87:80] : _GEN_1367; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1512 = 8'h47 == _T_22 ? io_in_bits[87:80] : _GEN_1368; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1513 = 8'h48 == _T_22 ? io_in_bits[87:80] : _GEN_1369; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1514 = 8'h49 == _T_22 ? io_in_bits[87:80] : _GEN_1370; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1515 = 8'h4a == _T_22 ? io_in_bits[87:80] : _GEN_1371; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1516 = 8'h4b == _T_22 ? io_in_bits[87:80] : _GEN_1372; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1517 = 8'h4c == _T_22 ? io_in_bits[87:80] : _GEN_1373; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1518 = 8'h4d == _T_22 ? io_in_bits[87:80] : _GEN_1374; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1519 = 8'h4e == _T_22 ? io_in_bits[87:80] : _GEN_1375; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1520 = 8'h4f == _T_22 ? io_in_bits[87:80] : _GEN_1376; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1521 = 8'h50 == _T_22 ? io_in_bits[87:80] : _GEN_1377; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1522 = 8'h51 == _T_22 ? io_in_bits[87:80] : _GEN_1378; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1523 = 8'h52 == _T_22 ? io_in_bits[87:80] : _GEN_1379; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1524 = 8'h53 == _T_22 ? io_in_bits[87:80] : _GEN_1380; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1525 = 8'h54 == _T_22 ? io_in_bits[87:80] : _GEN_1381; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1526 = 8'h55 == _T_22 ? io_in_bits[87:80] : _GEN_1382; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1527 = 8'h56 == _T_22 ? io_in_bits[87:80] : _GEN_1383; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1528 = 8'h57 == _T_22 ? io_in_bits[87:80] : _GEN_1384; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1529 = 8'h58 == _T_22 ? io_in_bits[87:80] : _GEN_1385; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1530 = 8'h59 == _T_22 ? io_in_bits[87:80] : _GEN_1386; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1531 = 8'h5a == _T_22 ? io_in_bits[87:80] : _GEN_1387; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1532 = 8'h5b == _T_22 ? io_in_bits[87:80] : _GEN_1388; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1533 = 8'h5c == _T_22 ? io_in_bits[87:80] : _GEN_1389; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1534 = 8'h5d == _T_22 ? io_in_bits[87:80] : _GEN_1390; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1535 = 8'h5e == _T_22 ? io_in_bits[87:80] : _GEN_1391; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1536 = 8'h5f == _T_22 ? io_in_bits[87:80] : _GEN_1392; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1537 = 8'h60 == _T_22 ? io_in_bits[87:80] : _GEN_1393; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1538 = 8'h61 == _T_22 ? io_in_bits[87:80] : _GEN_1394; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1539 = 8'h62 == _T_22 ? io_in_bits[87:80] : _GEN_1395; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1540 = 8'h63 == _T_22 ? io_in_bits[87:80] : _GEN_1396; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1541 = 8'h64 == _T_22 ? io_in_bits[87:80] : _GEN_1397; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1542 = 8'h65 == _T_22 ? io_in_bits[87:80] : _GEN_1398; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1543 = 8'h66 == _T_22 ? io_in_bits[87:80] : _GEN_1399; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1544 = 8'h67 == _T_22 ? io_in_bits[87:80] : _GEN_1400; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1545 = 8'h68 == _T_22 ? io_in_bits[87:80] : _GEN_1401; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1546 = 8'h69 == _T_22 ? io_in_bits[87:80] : _GEN_1402; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1547 = 8'h6a == _T_22 ? io_in_bits[87:80] : _GEN_1403; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1548 = 8'h6b == _T_22 ? io_in_bits[87:80] : _GEN_1404; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1549 = 8'h6c == _T_22 ? io_in_bits[87:80] : _GEN_1405; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1550 = 8'h6d == _T_22 ? io_in_bits[87:80] : _GEN_1406; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1551 = 8'h6e == _T_22 ? io_in_bits[87:80] : _GEN_1407; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1552 = 8'h6f == _T_22 ? io_in_bits[87:80] : _GEN_1408; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1553 = 8'h70 == _T_22 ? io_in_bits[87:80] : _GEN_1409; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1554 = 8'h71 == _T_22 ? io_in_bits[87:80] : _GEN_1410; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1555 = 8'h72 == _T_22 ? io_in_bits[87:80] : _GEN_1411; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1556 = 8'h73 == _T_22 ? io_in_bits[87:80] : _GEN_1412; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1557 = 8'h74 == _T_22 ? io_in_bits[87:80] : _GEN_1413; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1558 = 8'h75 == _T_22 ? io_in_bits[87:80] : _GEN_1414; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1559 = 8'h76 == _T_22 ? io_in_bits[87:80] : _GEN_1415; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1560 = 8'h77 == _T_22 ? io_in_bits[87:80] : _GEN_1416; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1561 = 8'h78 == _T_22 ? io_in_bits[87:80] : _GEN_1417; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1562 = 8'h79 == _T_22 ? io_in_bits[87:80] : _GEN_1418; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1563 = 8'h7a == _T_22 ? io_in_bits[87:80] : _GEN_1419; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1564 = 8'h7b == _T_22 ? io_in_bits[87:80] : _GEN_1420; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1565 = 8'h7c == _T_22 ? io_in_bits[87:80] : _GEN_1421; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1566 = 8'h7d == _T_22 ? io_in_bits[87:80] : _GEN_1422; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1567 = 8'h7e == _T_22 ? io_in_bits[87:80] : _GEN_1423; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1568 = 8'h7f == _T_22 ? io_in_bits[87:80] : _GEN_1424; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1569 = 8'h80 == _T_22 ? io_in_bits[87:80] : _GEN_1425; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1570 = 8'h81 == _T_22 ? io_in_bits[87:80] : _GEN_1426; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1571 = 8'h82 == _T_22 ? io_in_bits[87:80] : _GEN_1427; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1572 = 8'h83 == _T_22 ? io_in_bits[87:80] : _GEN_1428; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1573 = 8'h84 == _T_22 ? io_in_bits[87:80] : _GEN_1429; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1574 = 8'h85 == _T_22 ? io_in_bits[87:80] : _GEN_1430; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1575 = 8'h86 == _T_22 ? io_in_bits[87:80] : _GEN_1431; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1576 = 8'h87 == _T_22 ? io_in_bits[87:80] : _GEN_1432; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1577 = 8'h88 == _T_22 ? io_in_bits[87:80] : _GEN_1433; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1578 = 8'h89 == _T_22 ? io_in_bits[87:80] : _GEN_1434; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1579 = 8'h8a == _T_22 ? io_in_bits[87:80] : _GEN_1435; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1580 = 8'h8b == _T_22 ? io_in_bits[87:80] : _GEN_1436; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1581 = 8'h8c == _T_22 ? io_in_bits[87:80] : _GEN_1437; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1582 = 8'h8d == _T_22 ? io_in_bits[87:80] : _GEN_1438; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1583 = 8'h8e == _T_22 ? io_in_bits[87:80] : _GEN_1439; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1584 = 8'h8f == _T_22 ? io_in_bits[87:80] : _GEN_1440; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_24 = enqPtr + 8'hb; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_1585 = 8'h0 == _T_24 ? io_in_bits[95:88] : _GEN_1441; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1586 = 8'h1 == _T_24 ? io_in_bits[95:88] : _GEN_1442; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1587 = 8'h2 == _T_24 ? io_in_bits[95:88] : _GEN_1443; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1588 = 8'h3 == _T_24 ? io_in_bits[95:88] : _GEN_1444; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1589 = 8'h4 == _T_24 ? io_in_bits[95:88] : _GEN_1445; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1590 = 8'h5 == _T_24 ? io_in_bits[95:88] : _GEN_1446; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1591 = 8'h6 == _T_24 ? io_in_bits[95:88] : _GEN_1447; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1592 = 8'h7 == _T_24 ? io_in_bits[95:88] : _GEN_1448; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1593 = 8'h8 == _T_24 ? io_in_bits[95:88] : _GEN_1449; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1594 = 8'h9 == _T_24 ? io_in_bits[95:88] : _GEN_1450; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1595 = 8'ha == _T_24 ? io_in_bits[95:88] : _GEN_1451; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1596 = 8'hb == _T_24 ? io_in_bits[95:88] : _GEN_1452; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1597 = 8'hc == _T_24 ? io_in_bits[95:88] : _GEN_1453; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1598 = 8'hd == _T_24 ? io_in_bits[95:88] : _GEN_1454; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1599 = 8'he == _T_24 ? io_in_bits[95:88] : _GEN_1455; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1600 = 8'hf == _T_24 ? io_in_bits[95:88] : _GEN_1456; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1601 = 8'h10 == _T_24 ? io_in_bits[95:88] : _GEN_1457; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1602 = 8'h11 == _T_24 ? io_in_bits[95:88] : _GEN_1458; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1603 = 8'h12 == _T_24 ? io_in_bits[95:88] : _GEN_1459; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1604 = 8'h13 == _T_24 ? io_in_bits[95:88] : _GEN_1460; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1605 = 8'h14 == _T_24 ? io_in_bits[95:88] : _GEN_1461; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1606 = 8'h15 == _T_24 ? io_in_bits[95:88] : _GEN_1462; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1607 = 8'h16 == _T_24 ? io_in_bits[95:88] : _GEN_1463; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1608 = 8'h17 == _T_24 ? io_in_bits[95:88] : _GEN_1464; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1609 = 8'h18 == _T_24 ? io_in_bits[95:88] : _GEN_1465; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1610 = 8'h19 == _T_24 ? io_in_bits[95:88] : _GEN_1466; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1611 = 8'h1a == _T_24 ? io_in_bits[95:88] : _GEN_1467; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1612 = 8'h1b == _T_24 ? io_in_bits[95:88] : _GEN_1468; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1613 = 8'h1c == _T_24 ? io_in_bits[95:88] : _GEN_1469; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1614 = 8'h1d == _T_24 ? io_in_bits[95:88] : _GEN_1470; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1615 = 8'h1e == _T_24 ? io_in_bits[95:88] : _GEN_1471; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1616 = 8'h1f == _T_24 ? io_in_bits[95:88] : _GEN_1472; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1617 = 8'h20 == _T_24 ? io_in_bits[95:88] : _GEN_1473; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1618 = 8'h21 == _T_24 ? io_in_bits[95:88] : _GEN_1474; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1619 = 8'h22 == _T_24 ? io_in_bits[95:88] : _GEN_1475; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1620 = 8'h23 == _T_24 ? io_in_bits[95:88] : _GEN_1476; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1621 = 8'h24 == _T_24 ? io_in_bits[95:88] : _GEN_1477; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1622 = 8'h25 == _T_24 ? io_in_bits[95:88] : _GEN_1478; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1623 = 8'h26 == _T_24 ? io_in_bits[95:88] : _GEN_1479; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1624 = 8'h27 == _T_24 ? io_in_bits[95:88] : _GEN_1480; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1625 = 8'h28 == _T_24 ? io_in_bits[95:88] : _GEN_1481; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1626 = 8'h29 == _T_24 ? io_in_bits[95:88] : _GEN_1482; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1627 = 8'h2a == _T_24 ? io_in_bits[95:88] : _GEN_1483; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1628 = 8'h2b == _T_24 ? io_in_bits[95:88] : _GEN_1484; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1629 = 8'h2c == _T_24 ? io_in_bits[95:88] : _GEN_1485; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1630 = 8'h2d == _T_24 ? io_in_bits[95:88] : _GEN_1486; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1631 = 8'h2e == _T_24 ? io_in_bits[95:88] : _GEN_1487; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1632 = 8'h2f == _T_24 ? io_in_bits[95:88] : _GEN_1488; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1633 = 8'h30 == _T_24 ? io_in_bits[95:88] : _GEN_1489; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1634 = 8'h31 == _T_24 ? io_in_bits[95:88] : _GEN_1490; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1635 = 8'h32 == _T_24 ? io_in_bits[95:88] : _GEN_1491; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1636 = 8'h33 == _T_24 ? io_in_bits[95:88] : _GEN_1492; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1637 = 8'h34 == _T_24 ? io_in_bits[95:88] : _GEN_1493; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1638 = 8'h35 == _T_24 ? io_in_bits[95:88] : _GEN_1494; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1639 = 8'h36 == _T_24 ? io_in_bits[95:88] : _GEN_1495; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1640 = 8'h37 == _T_24 ? io_in_bits[95:88] : _GEN_1496; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1641 = 8'h38 == _T_24 ? io_in_bits[95:88] : _GEN_1497; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1642 = 8'h39 == _T_24 ? io_in_bits[95:88] : _GEN_1498; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1643 = 8'h3a == _T_24 ? io_in_bits[95:88] : _GEN_1499; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1644 = 8'h3b == _T_24 ? io_in_bits[95:88] : _GEN_1500; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1645 = 8'h3c == _T_24 ? io_in_bits[95:88] : _GEN_1501; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1646 = 8'h3d == _T_24 ? io_in_bits[95:88] : _GEN_1502; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1647 = 8'h3e == _T_24 ? io_in_bits[95:88] : _GEN_1503; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1648 = 8'h3f == _T_24 ? io_in_bits[95:88] : _GEN_1504; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1649 = 8'h40 == _T_24 ? io_in_bits[95:88] : _GEN_1505; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1650 = 8'h41 == _T_24 ? io_in_bits[95:88] : _GEN_1506; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1651 = 8'h42 == _T_24 ? io_in_bits[95:88] : _GEN_1507; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1652 = 8'h43 == _T_24 ? io_in_bits[95:88] : _GEN_1508; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1653 = 8'h44 == _T_24 ? io_in_bits[95:88] : _GEN_1509; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1654 = 8'h45 == _T_24 ? io_in_bits[95:88] : _GEN_1510; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1655 = 8'h46 == _T_24 ? io_in_bits[95:88] : _GEN_1511; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1656 = 8'h47 == _T_24 ? io_in_bits[95:88] : _GEN_1512; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1657 = 8'h48 == _T_24 ? io_in_bits[95:88] : _GEN_1513; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1658 = 8'h49 == _T_24 ? io_in_bits[95:88] : _GEN_1514; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1659 = 8'h4a == _T_24 ? io_in_bits[95:88] : _GEN_1515; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1660 = 8'h4b == _T_24 ? io_in_bits[95:88] : _GEN_1516; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1661 = 8'h4c == _T_24 ? io_in_bits[95:88] : _GEN_1517; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1662 = 8'h4d == _T_24 ? io_in_bits[95:88] : _GEN_1518; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1663 = 8'h4e == _T_24 ? io_in_bits[95:88] : _GEN_1519; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1664 = 8'h4f == _T_24 ? io_in_bits[95:88] : _GEN_1520; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1665 = 8'h50 == _T_24 ? io_in_bits[95:88] : _GEN_1521; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1666 = 8'h51 == _T_24 ? io_in_bits[95:88] : _GEN_1522; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1667 = 8'h52 == _T_24 ? io_in_bits[95:88] : _GEN_1523; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1668 = 8'h53 == _T_24 ? io_in_bits[95:88] : _GEN_1524; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1669 = 8'h54 == _T_24 ? io_in_bits[95:88] : _GEN_1525; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1670 = 8'h55 == _T_24 ? io_in_bits[95:88] : _GEN_1526; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1671 = 8'h56 == _T_24 ? io_in_bits[95:88] : _GEN_1527; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1672 = 8'h57 == _T_24 ? io_in_bits[95:88] : _GEN_1528; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1673 = 8'h58 == _T_24 ? io_in_bits[95:88] : _GEN_1529; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1674 = 8'h59 == _T_24 ? io_in_bits[95:88] : _GEN_1530; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1675 = 8'h5a == _T_24 ? io_in_bits[95:88] : _GEN_1531; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1676 = 8'h5b == _T_24 ? io_in_bits[95:88] : _GEN_1532; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1677 = 8'h5c == _T_24 ? io_in_bits[95:88] : _GEN_1533; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1678 = 8'h5d == _T_24 ? io_in_bits[95:88] : _GEN_1534; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1679 = 8'h5e == _T_24 ? io_in_bits[95:88] : _GEN_1535; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1680 = 8'h5f == _T_24 ? io_in_bits[95:88] : _GEN_1536; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1681 = 8'h60 == _T_24 ? io_in_bits[95:88] : _GEN_1537; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1682 = 8'h61 == _T_24 ? io_in_bits[95:88] : _GEN_1538; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1683 = 8'h62 == _T_24 ? io_in_bits[95:88] : _GEN_1539; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1684 = 8'h63 == _T_24 ? io_in_bits[95:88] : _GEN_1540; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1685 = 8'h64 == _T_24 ? io_in_bits[95:88] : _GEN_1541; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1686 = 8'h65 == _T_24 ? io_in_bits[95:88] : _GEN_1542; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1687 = 8'h66 == _T_24 ? io_in_bits[95:88] : _GEN_1543; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1688 = 8'h67 == _T_24 ? io_in_bits[95:88] : _GEN_1544; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1689 = 8'h68 == _T_24 ? io_in_bits[95:88] : _GEN_1545; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1690 = 8'h69 == _T_24 ? io_in_bits[95:88] : _GEN_1546; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1691 = 8'h6a == _T_24 ? io_in_bits[95:88] : _GEN_1547; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1692 = 8'h6b == _T_24 ? io_in_bits[95:88] : _GEN_1548; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1693 = 8'h6c == _T_24 ? io_in_bits[95:88] : _GEN_1549; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1694 = 8'h6d == _T_24 ? io_in_bits[95:88] : _GEN_1550; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1695 = 8'h6e == _T_24 ? io_in_bits[95:88] : _GEN_1551; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1696 = 8'h6f == _T_24 ? io_in_bits[95:88] : _GEN_1552; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1697 = 8'h70 == _T_24 ? io_in_bits[95:88] : _GEN_1553; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1698 = 8'h71 == _T_24 ? io_in_bits[95:88] : _GEN_1554; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1699 = 8'h72 == _T_24 ? io_in_bits[95:88] : _GEN_1555; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1700 = 8'h73 == _T_24 ? io_in_bits[95:88] : _GEN_1556; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1701 = 8'h74 == _T_24 ? io_in_bits[95:88] : _GEN_1557; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1702 = 8'h75 == _T_24 ? io_in_bits[95:88] : _GEN_1558; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1703 = 8'h76 == _T_24 ? io_in_bits[95:88] : _GEN_1559; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1704 = 8'h77 == _T_24 ? io_in_bits[95:88] : _GEN_1560; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1705 = 8'h78 == _T_24 ? io_in_bits[95:88] : _GEN_1561; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1706 = 8'h79 == _T_24 ? io_in_bits[95:88] : _GEN_1562; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1707 = 8'h7a == _T_24 ? io_in_bits[95:88] : _GEN_1563; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1708 = 8'h7b == _T_24 ? io_in_bits[95:88] : _GEN_1564; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1709 = 8'h7c == _T_24 ? io_in_bits[95:88] : _GEN_1565; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1710 = 8'h7d == _T_24 ? io_in_bits[95:88] : _GEN_1566; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1711 = 8'h7e == _T_24 ? io_in_bits[95:88] : _GEN_1567; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1712 = 8'h7f == _T_24 ? io_in_bits[95:88] : _GEN_1568; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1713 = 8'h80 == _T_24 ? io_in_bits[95:88] : _GEN_1569; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1714 = 8'h81 == _T_24 ? io_in_bits[95:88] : _GEN_1570; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1715 = 8'h82 == _T_24 ? io_in_bits[95:88] : _GEN_1571; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1716 = 8'h83 == _T_24 ? io_in_bits[95:88] : _GEN_1572; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1717 = 8'h84 == _T_24 ? io_in_bits[95:88] : _GEN_1573; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1718 = 8'h85 == _T_24 ? io_in_bits[95:88] : _GEN_1574; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1719 = 8'h86 == _T_24 ? io_in_bits[95:88] : _GEN_1575; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1720 = 8'h87 == _T_24 ? io_in_bits[95:88] : _GEN_1576; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1721 = 8'h88 == _T_24 ? io_in_bits[95:88] : _GEN_1577; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1722 = 8'h89 == _T_24 ? io_in_bits[95:88] : _GEN_1578; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1723 = 8'h8a == _T_24 ? io_in_bits[95:88] : _GEN_1579; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1724 = 8'h8b == _T_24 ? io_in_bits[95:88] : _GEN_1580; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1725 = 8'h8c == _T_24 ? io_in_bits[95:88] : _GEN_1581; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1726 = 8'h8d == _T_24 ? io_in_bits[95:88] : _GEN_1582; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1727 = 8'h8e == _T_24 ? io_in_bits[95:88] : _GEN_1583; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1728 = 8'h8f == _T_24 ? io_in_bits[95:88] : _GEN_1584; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_26 = enqPtr + 8'hc; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_1729 = 8'h0 == _T_26 ? io_in_bits[103:96] : _GEN_1585; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1730 = 8'h1 == _T_26 ? io_in_bits[103:96] : _GEN_1586; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1731 = 8'h2 == _T_26 ? io_in_bits[103:96] : _GEN_1587; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1732 = 8'h3 == _T_26 ? io_in_bits[103:96] : _GEN_1588; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1733 = 8'h4 == _T_26 ? io_in_bits[103:96] : _GEN_1589; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1734 = 8'h5 == _T_26 ? io_in_bits[103:96] : _GEN_1590; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1735 = 8'h6 == _T_26 ? io_in_bits[103:96] : _GEN_1591; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1736 = 8'h7 == _T_26 ? io_in_bits[103:96] : _GEN_1592; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1737 = 8'h8 == _T_26 ? io_in_bits[103:96] : _GEN_1593; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1738 = 8'h9 == _T_26 ? io_in_bits[103:96] : _GEN_1594; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1739 = 8'ha == _T_26 ? io_in_bits[103:96] : _GEN_1595; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1740 = 8'hb == _T_26 ? io_in_bits[103:96] : _GEN_1596; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1741 = 8'hc == _T_26 ? io_in_bits[103:96] : _GEN_1597; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1742 = 8'hd == _T_26 ? io_in_bits[103:96] : _GEN_1598; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1743 = 8'he == _T_26 ? io_in_bits[103:96] : _GEN_1599; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1744 = 8'hf == _T_26 ? io_in_bits[103:96] : _GEN_1600; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1745 = 8'h10 == _T_26 ? io_in_bits[103:96] : _GEN_1601; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1746 = 8'h11 == _T_26 ? io_in_bits[103:96] : _GEN_1602; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1747 = 8'h12 == _T_26 ? io_in_bits[103:96] : _GEN_1603; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1748 = 8'h13 == _T_26 ? io_in_bits[103:96] : _GEN_1604; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1749 = 8'h14 == _T_26 ? io_in_bits[103:96] : _GEN_1605; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1750 = 8'h15 == _T_26 ? io_in_bits[103:96] : _GEN_1606; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1751 = 8'h16 == _T_26 ? io_in_bits[103:96] : _GEN_1607; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1752 = 8'h17 == _T_26 ? io_in_bits[103:96] : _GEN_1608; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1753 = 8'h18 == _T_26 ? io_in_bits[103:96] : _GEN_1609; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1754 = 8'h19 == _T_26 ? io_in_bits[103:96] : _GEN_1610; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1755 = 8'h1a == _T_26 ? io_in_bits[103:96] : _GEN_1611; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1756 = 8'h1b == _T_26 ? io_in_bits[103:96] : _GEN_1612; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1757 = 8'h1c == _T_26 ? io_in_bits[103:96] : _GEN_1613; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1758 = 8'h1d == _T_26 ? io_in_bits[103:96] : _GEN_1614; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1759 = 8'h1e == _T_26 ? io_in_bits[103:96] : _GEN_1615; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1760 = 8'h1f == _T_26 ? io_in_bits[103:96] : _GEN_1616; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1761 = 8'h20 == _T_26 ? io_in_bits[103:96] : _GEN_1617; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1762 = 8'h21 == _T_26 ? io_in_bits[103:96] : _GEN_1618; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1763 = 8'h22 == _T_26 ? io_in_bits[103:96] : _GEN_1619; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1764 = 8'h23 == _T_26 ? io_in_bits[103:96] : _GEN_1620; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1765 = 8'h24 == _T_26 ? io_in_bits[103:96] : _GEN_1621; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1766 = 8'h25 == _T_26 ? io_in_bits[103:96] : _GEN_1622; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1767 = 8'h26 == _T_26 ? io_in_bits[103:96] : _GEN_1623; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1768 = 8'h27 == _T_26 ? io_in_bits[103:96] : _GEN_1624; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1769 = 8'h28 == _T_26 ? io_in_bits[103:96] : _GEN_1625; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1770 = 8'h29 == _T_26 ? io_in_bits[103:96] : _GEN_1626; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1771 = 8'h2a == _T_26 ? io_in_bits[103:96] : _GEN_1627; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1772 = 8'h2b == _T_26 ? io_in_bits[103:96] : _GEN_1628; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1773 = 8'h2c == _T_26 ? io_in_bits[103:96] : _GEN_1629; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1774 = 8'h2d == _T_26 ? io_in_bits[103:96] : _GEN_1630; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1775 = 8'h2e == _T_26 ? io_in_bits[103:96] : _GEN_1631; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1776 = 8'h2f == _T_26 ? io_in_bits[103:96] : _GEN_1632; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1777 = 8'h30 == _T_26 ? io_in_bits[103:96] : _GEN_1633; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1778 = 8'h31 == _T_26 ? io_in_bits[103:96] : _GEN_1634; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1779 = 8'h32 == _T_26 ? io_in_bits[103:96] : _GEN_1635; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1780 = 8'h33 == _T_26 ? io_in_bits[103:96] : _GEN_1636; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1781 = 8'h34 == _T_26 ? io_in_bits[103:96] : _GEN_1637; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1782 = 8'h35 == _T_26 ? io_in_bits[103:96] : _GEN_1638; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1783 = 8'h36 == _T_26 ? io_in_bits[103:96] : _GEN_1639; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1784 = 8'h37 == _T_26 ? io_in_bits[103:96] : _GEN_1640; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1785 = 8'h38 == _T_26 ? io_in_bits[103:96] : _GEN_1641; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1786 = 8'h39 == _T_26 ? io_in_bits[103:96] : _GEN_1642; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1787 = 8'h3a == _T_26 ? io_in_bits[103:96] : _GEN_1643; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1788 = 8'h3b == _T_26 ? io_in_bits[103:96] : _GEN_1644; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1789 = 8'h3c == _T_26 ? io_in_bits[103:96] : _GEN_1645; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1790 = 8'h3d == _T_26 ? io_in_bits[103:96] : _GEN_1646; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1791 = 8'h3e == _T_26 ? io_in_bits[103:96] : _GEN_1647; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1792 = 8'h3f == _T_26 ? io_in_bits[103:96] : _GEN_1648; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1793 = 8'h40 == _T_26 ? io_in_bits[103:96] : _GEN_1649; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1794 = 8'h41 == _T_26 ? io_in_bits[103:96] : _GEN_1650; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1795 = 8'h42 == _T_26 ? io_in_bits[103:96] : _GEN_1651; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1796 = 8'h43 == _T_26 ? io_in_bits[103:96] : _GEN_1652; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1797 = 8'h44 == _T_26 ? io_in_bits[103:96] : _GEN_1653; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1798 = 8'h45 == _T_26 ? io_in_bits[103:96] : _GEN_1654; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1799 = 8'h46 == _T_26 ? io_in_bits[103:96] : _GEN_1655; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1800 = 8'h47 == _T_26 ? io_in_bits[103:96] : _GEN_1656; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1801 = 8'h48 == _T_26 ? io_in_bits[103:96] : _GEN_1657; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1802 = 8'h49 == _T_26 ? io_in_bits[103:96] : _GEN_1658; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1803 = 8'h4a == _T_26 ? io_in_bits[103:96] : _GEN_1659; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1804 = 8'h4b == _T_26 ? io_in_bits[103:96] : _GEN_1660; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1805 = 8'h4c == _T_26 ? io_in_bits[103:96] : _GEN_1661; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1806 = 8'h4d == _T_26 ? io_in_bits[103:96] : _GEN_1662; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1807 = 8'h4e == _T_26 ? io_in_bits[103:96] : _GEN_1663; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1808 = 8'h4f == _T_26 ? io_in_bits[103:96] : _GEN_1664; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1809 = 8'h50 == _T_26 ? io_in_bits[103:96] : _GEN_1665; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1810 = 8'h51 == _T_26 ? io_in_bits[103:96] : _GEN_1666; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1811 = 8'h52 == _T_26 ? io_in_bits[103:96] : _GEN_1667; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1812 = 8'h53 == _T_26 ? io_in_bits[103:96] : _GEN_1668; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1813 = 8'h54 == _T_26 ? io_in_bits[103:96] : _GEN_1669; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1814 = 8'h55 == _T_26 ? io_in_bits[103:96] : _GEN_1670; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1815 = 8'h56 == _T_26 ? io_in_bits[103:96] : _GEN_1671; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1816 = 8'h57 == _T_26 ? io_in_bits[103:96] : _GEN_1672; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1817 = 8'h58 == _T_26 ? io_in_bits[103:96] : _GEN_1673; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1818 = 8'h59 == _T_26 ? io_in_bits[103:96] : _GEN_1674; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1819 = 8'h5a == _T_26 ? io_in_bits[103:96] : _GEN_1675; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1820 = 8'h5b == _T_26 ? io_in_bits[103:96] : _GEN_1676; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1821 = 8'h5c == _T_26 ? io_in_bits[103:96] : _GEN_1677; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1822 = 8'h5d == _T_26 ? io_in_bits[103:96] : _GEN_1678; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1823 = 8'h5e == _T_26 ? io_in_bits[103:96] : _GEN_1679; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1824 = 8'h5f == _T_26 ? io_in_bits[103:96] : _GEN_1680; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1825 = 8'h60 == _T_26 ? io_in_bits[103:96] : _GEN_1681; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1826 = 8'h61 == _T_26 ? io_in_bits[103:96] : _GEN_1682; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1827 = 8'h62 == _T_26 ? io_in_bits[103:96] : _GEN_1683; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1828 = 8'h63 == _T_26 ? io_in_bits[103:96] : _GEN_1684; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1829 = 8'h64 == _T_26 ? io_in_bits[103:96] : _GEN_1685; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1830 = 8'h65 == _T_26 ? io_in_bits[103:96] : _GEN_1686; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1831 = 8'h66 == _T_26 ? io_in_bits[103:96] : _GEN_1687; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1832 = 8'h67 == _T_26 ? io_in_bits[103:96] : _GEN_1688; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1833 = 8'h68 == _T_26 ? io_in_bits[103:96] : _GEN_1689; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1834 = 8'h69 == _T_26 ? io_in_bits[103:96] : _GEN_1690; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1835 = 8'h6a == _T_26 ? io_in_bits[103:96] : _GEN_1691; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1836 = 8'h6b == _T_26 ? io_in_bits[103:96] : _GEN_1692; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1837 = 8'h6c == _T_26 ? io_in_bits[103:96] : _GEN_1693; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1838 = 8'h6d == _T_26 ? io_in_bits[103:96] : _GEN_1694; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1839 = 8'h6e == _T_26 ? io_in_bits[103:96] : _GEN_1695; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1840 = 8'h6f == _T_26 ? io_in_bits[103:96] : _GEN_1696; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1841 = 8'h70 == _T_26 ? io_in_bits[103:96] : _GEN_1697; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1842 = 8'h71 == _T_26 ? io_in_bits[103:96] : _GEN_1698; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1843 = 8'h72 == _T_26 ? io_in_bits[103:96] : _GEN_1699; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1844 = 8'h73 == _T_26 ? io_in_bits[103:96] : _GEN_1700; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1845 = 8'h74 == _T_26 ? io_in_bits[103:96] : _GEN_1701; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1846 = 8'h75 == _T_26 ? io_in_bits[103:96] : _GEN_1702; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1847 = 8'h76 == _T_26 ? io_in_bits[103:96] : _GEN_1703; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1848 = 8'h77 == _T_26 ? io_in_bits[103:96] : _GEN_1704; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1849 = 8'h78 == _T_26 ? io_in_bits[103:96] : _GEN_1705; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1850 = 8'h79 == _T_26 ? io_in_bits[103:96] : _GEN_1706; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1851 = 8'h7a == _T_26 ? io_in_bits[103:96] : _GEN_1707; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1852 = 8'h7b == _T_26 ? io_in_bits[103:96] : _GEN_1708; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1853 = 8'h7c == _T_26 ? io_in_bits[103:96] : _GEN_1709; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1854 = 8'h7d == _T_26 ? io_in_bits[103:96] : _GEN_1710; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1855 = 8'h7e == _T_26 ? io_in_bits[103:96] : _GEN_1711; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1856 = 8'h7f == _T_26 ? io_in_bits[103:96] : _GEN_1712; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1857 = 8'h80 == _T_26 ? io_in_bits[103:96] : _GEN_1713; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1858 = 8'h81 == _T_26 ? io_in_bits[103:96] : _GEN_1714; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1859 = 8'h82 == _T_26 ? io_in_bits[103:96] : _GEN_1715; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1860 = 8'h83 == _T_26 ? io_in_bits[103:96] : _GEN_1716; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1861 = 8'h84 == _T_26 ? io_in_bits[103:96] : _GEN_1717; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1862 = 8'h85 == _T_26 ? io_in_bits[103:96] : _GEN_1718; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1863 = 8'h86 == _T_26 ? io_in_bits[103:96] : _GEN_1719; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1864 = 8'h87 == _T_26 ? io_in_bits[103:96] : _GEN_1720; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1865 = 8'h88 == _T_26 ? io_in_bits[103:96] : _GEN_1721; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1866 = 8'h89 == _T_26 ? io_in_bits[103:96] : _GEN_1722; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1867 = 8'h8a == _T_26 ? io_in_bits[103:96] : _GEN_1723; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1868 = 8'h8b == _T_26 ? io_in_bits[103:96] : _GEN_1724; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1869 = 8'h8c == _T_26 ? io_in_bits[103:96] : _GEN_1725; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1870 = 8'h8d == _T_26 ? io_in_bits[103:96] : _GEN_1726; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1871 = 8'h8e == _T_26 ? io_in_bits[103:96] : _GEN_1727; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1872 = 8'h8f == _T_26 ? io_in_bits[103:96] : _GEN_1728; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_28 = enqPtr + 8'hd; // @[WidthConverter.scala 67:20]
  wire [7:0] _GEN_1873 = 8'h0 == _T_28 ? io_in_bits[111:104] : _GEN_1729; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1874 = 8'h1 == _T_28 ? io_in_bits[111:104] : _GEN_1730; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1875 = 8'h2 == _T_28 ? io_in_bits[111:104] : _GEN_1731; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1876 = 8'h3 == _T_28 ? io_in_bits[111:104] : _GEN_1732; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1877 = 8'h4 == _T_28 ? io_in_bits[111:104] : _GEN_1733; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1878 = 8'h5 == _T_28 ? io_in_bits[111:104] : _GEN_1734; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1879 = 8'h6 == _T_28 ? io_in_bits[111:104] : _GEN_1735; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1880 = 8'h7 == _T_28 ? io_in_bits[111:104] : _GEN_1736; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1881 = 8'h8 == _T_28 ? io_in_bits[111:104] : _GEN_1737; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1882 = 8'h9 == _T_28 ? io_in_bits[111:104] : _GEN_1738; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1883 = 8'ha == _T_28 ? io_in_bits[111:104] : _GEN_1739; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1884 = 8'hb == _T_28 ? io_in_bits[111:104] : _GEN_1740; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1885 = 8'hc == _T_28 ? io_in_bits[111:104] : _GEN_1741; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1886 = 8'hd == _T_28 ? io_in_bits[111:104] : _GEN_1742; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1887 = 8'he == _T_28 ? io_in_bits[111:104] : _GEN_1743; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1888 = 8'hf == _T_28 ? io_in_bits[111:104] : _GEN_1744; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1889 = 8'h10 == _T_28 ? io_in_bits[111:104] : _GEN_1745; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1890 = 8'h11 == _T_28 ? io_in_bits[111:104] : _GEN_1746; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1891 = 8'h12 == _T_28 ? io_in_bits[111:104] : _GEN_1747; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1892 = 8'h13 == _T_28 ? io_in_bits[111:104] : _GEN_1748; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1893 = 8'h14 == _T_28 ? io_in_bits[111:104] : _GEN_1749; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1894 = 8'h15 == _T_28 ? io_in_bits[111:104] : _GEN_1750; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1895 = 8'h16 == _T_28 ? io_in_bits[111:104] : _GEN_1751; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1896 = 8'h17 == _T_28 ? io_in_bits[111:104] : _GEN_1752; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1897 = 8'h18 == _T_28 ? io_in_bits[111:104] : _GEN_1753; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1898 = 8'h19 == _T_28 ? io_in_bits[111:104] : _GEN_1754; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1899 = 8'h1a == _T_28 ? io_in_bits[111:104] : _GEN_1755; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1900 = 8'h1b == _T_28 ? io_in_bits[111:104] : _GEN_1756; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1901 = 8'h1c == _T_28 ? io_in_bits[111:104] : _GEN_1757; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1902 = 8'h1d == _T_28 ? io_in_bits[111:104] : _GEN_1758; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1903 = 8'h1e == _T_28 ? io_in_bits[111:104] : _GEN_1759; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1904 = 8'h1f == _T_28 ? io_in_bits[111:104] : _GEN_1760; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1905 = 8'h20 == _T_28 ? io_in_bits[111:104] : _GEN_1761; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1906 = 8'h21 == _T_28 ? io_in_bits[111:104] : _GEN_1762; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1907 = 8'h22 == _T_28 ? io_in_bits[111:104] : _GEN_1763; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1908 = 8'h23 == _T_28 ? io_in_bits[111:104] : _GEN_1764; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1909 = 8'h24 == _T_28 ? io_in_bits[111:104] : _GEN_1765; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1910 = 8'h25 == _T_28 ? io_in_bits[111:104] : _GEN_1766; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1911 = 8'h26 == _T_28 ? io_in_bits[111:104] : _GEN_1767; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1912 = 8'h27 == _T_28 ? io_in_bits[111:104] : _GEN_1768; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1913 = 8'h28 == _T_28 ? io_in_bits[111:104] : _GEN_1769; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1914 = 8'h29 == _T_28 ? io_in_bits[111:104] : _GEN_1770; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1915 = 8'h2a == _T_28 ? io_in_bits[111:104] : _GEN_1771; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1916 = 8'h2b == _T_28 ? io_in_bits[111:104] : _GEN_1772; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1917 = 8'h2c == _T_28 ? io_in_bits[111:104] : _GEN_1773; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1918 = 8'h2d == _T_28 ? io_in_bits[111:104] : _GEN_1774; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1919 = 8'h2e == _T_28 ? io_in_bits[111:104] : _GEN_1775; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1920 = 8'h2f == _T_28 ? io_in_bits[111:104] : _GEN_1776; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1921 = 8'h30 == _T_28 ? io_in_bits[111:104] : _GEN_1777; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1922 = 8'h31 == _T_28 ? io_in_bits[111:104] : _GEN_1778; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1923 = 8'h32 == _T_28 ? io_in_bits[111:104] : _GEN_1779; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1924 = 8'h33 == _T_28 ? io_in_bits[111:104] : _GEN_1780; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1925 = 8'h34 == _T_28 ? io_in_bits[111:104] : _GEN_1781; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1926 = 8'h35 == _T_28 ? io_in_bits[111:104] : _GEN_1782; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1927 = 8'h36 == _T_28 ? io_in_bits[111:104] : _GEN_1783; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1928 = 8'h37 == _T_28 ? io_in_bits[111:104] : _GEN_1784; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1929 = 8'h38 == _T_28 ? io_in_bits[111:104] : _GEN_1785; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1930 = 8'h39 == _T_28 ? io_in_bits[111:104] : _GEN_1786; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1931 = 8'h3a == _T_28 ? io_in_bits[111:104] : _GEN_1787; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1932 = 8'h3b == _T_28 ? io_in_bits[111:104] : _GEN_1788; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1933 = 8'h3c == _T_28 ? io_in_bits[111:104] : _GEN_1789; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1934 = 8'h3d == _T_28 ? io_in_bits[111:104] : _GEN_1790; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1935 = 8'h3e == _T_28 ? io_in_bits[111:104] : _GEN_1791; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1936 = 8'h3f == _T_28 ? io_in_bits[111:104] : _GEN_1792; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1937 = 8'h40 == _T_28 ? io_in_bits[111:104] : _GEN_1793; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1938 = 8'h41 == _T_28 ? io_in_bits[111:104] : _GEN_1794; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1939 = 8'h42 == _T_28 ? io_in_bits[111:104] : _GEN_1795; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1940 = 8'h43 == _T_28 ? io_in_bits[111:104] : _GEN_1796; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1941 = 8'h44 == _T_28 ? io_in_bits[111:104] : _GEN_1797; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1942 = 8'h45 == _T_28 ? io_in_bits[111:104] : _GEN_1798; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1943 = 8'h46 == _T_28 ? io_in_bits[111:104] : _GEN_1799; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1944 = 8'h47 == _T_28 ? io_in_bits[111:104] : _GEN_1800; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1945 = 8'h48 == _T_28 ? io_in_bits[111:104] : _GEN_1801; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1946 = 8'h49 == _T_28 ? io_in_bits[111:104] : _GEN_1802; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1947 = 8'h4a == _T_28 ? io_in_bits[111:104] : _GEN_1803; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1948 = 8'h4b == _T_28 ? io_in_bits[111:104] : _GEN_1804; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1949 = 8'h4c == _T_28 ? io_in_bits[111:104] : _GEN_1805; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1950 = 8'h4d == _T_28 ? io_in_bits[111:104] : _GEN_1806; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1951 = 8'h4e == _T_28 ? io_in_bits[111:104] : _GEN_1807; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1952 = 8'h4f == _T_28 ? io_in_bits[111:104] : _GEN_1808; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1953 = 8'h50 == _T_28 ? io_in_bits[111:104] : _GEN_1809; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1954 = 8'h51 == _T_28 ? io_in_bits[111:104] : _GEN_1810; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1955 = 8'h52 == _T_28 ? io_in_bits[111:104] : _GEN_1811; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1956 = 8'h53 == _T_28 ? io_in_bits[111:104] : _GEN_1812; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1957 = 8'h54 == _T_28 ? io_in_bits[111:104] : _GEN_1813; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1958 = 8'h55 == _T_28 ? io_in_bits[111:104] : _GEN_1814; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1959 = 8'h56 == _T_28 ? io_in_bits[111:104] : _GEN_1815; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1960 = 8'h57 == _T_28 ? io_in_bits[111:104] : _GEN_1816; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1961 = 8'h58 == _T_28 ? io_in_bits[111:104] : _GEN_1817; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1962 = 8'h59 == _T_28 ? io_in_bits[111:104] : _GEN_1818; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1963 = 8'h5a == _T_28 ? io_in_bits[111:104] : _GEN_1819; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1964 = 8'h5b == _T_28 ? io_in_bits[111:104] : _GEN_1820; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1965 = 8'h5c == _T_28 ? io_in_bits[111:104] : _GEN_1821; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1966 = 8'h5d == _T_28 ? io_in_bits[111:104] : _GEN_1822; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1967 = 8'h5e == _T_28 ? io_in_bits[111:104] : _GEN_1823; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1968 = 8'h5f == _T_28 ? io_in_bits[111:104] : _GEN_1824; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1969 = 8'h60 == _T_28 ? io_in_bits[111:104] : _GEN_1825; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1970 = 8'h61 == _T_28 ? io_in_bits[111:104] : _GEN_1826; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1971 = 8'h62 == _T_28 ? io_in_bits[111:104] : _GEN_1827; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1972 = 8'h63 == _T_28 ? io_in_bits[111:104] : _GEN_1828; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1973 = 8'h64 == _T_28 ? io_in_bits[111:104] : _GEN_1829; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1974 = 8'h65 == _T_28 ? io_in_bits[111:104] : _GEN_1830; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1975 = 8'h66 == _T_28 ? io_in_bits[111:104] : _GEN_1831; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1976 = 8'h67 == _T_28 ? io_in_bits[111:104] : _GEN_1832; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1977 = 8'h68 == _T_28 ? io_in_bits[111:104] : _GEN_1833; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1978 = 8'h69 == _T_28 ? io_in_bits[111:104] : _GEN_1834; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1979 = 8'h6a == _T_28 ? io_in_bits[111:104] : _GEN_1835; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1980 = 8'h6b == _T_28 ? io_in_bits[111:104] : _GEN_1836; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1981 = 8'h6c == _T_28 ? io_in_bits[111:104] : _GEN_1837; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1982 = 8'h6d == _T_28 ? io_in_bits[111:104] : _GEN_1838; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1983 = 8'h6e == _T_28 ? io_in_bits[111:104] : _GEN_1839; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1984 = 8'h6f == _T_28 ? io_in_bits[111:104] : _GEN_1840; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1985 = 8'h70 == _T_28 ? io_in_bits[111:104] : _GEN_1841; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1986 = 8'h71 == _T_28 ? io_in_bits[111:104] : _GEN_1842; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1987 = 8'h72 == _T_28 ? io_in_bits[111:104] : _GEN_1843; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1988 = 8'h73 == _T_28 ? io_in_bits[111:104] : _GEN_1844; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1989 = 8'h74 == _T_28 ? io_in_bits[111:104] : _GEN_1845; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1990 = 8'h75 == _T_28 ? io_in_bits[111:104] : _GEN_1846; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1991 = 8'h76 == _T_28 ? io_in_bits[111:104] : _GEN_1847; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1992 = 8'h77 == _T_28 ? io_in_bits[111:104] : _GEN_1848; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1993 = 8'h78 == _T_28 ? io_in_bits[111:104] : _GEN_1849; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1994 = 8'h79 == _T_28 ? io_in_bits[111:104] : _GEN_1850; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1995 = 8'h7a == _T_28 ? io_in_bits[111:104] : _GEN_1851; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1996 = 8'h7b == _T_28 ? io_in_bits[111:104] : _GEN_1852; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1997 = 8'h7c == _T_28 ? io_in_bits[111:104] : _GEN_1853; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1998 = 8'h7d == _T_28 ? io_in_bits[111:104] : _GEN_1854; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_1999 = 8'h7e == _T_28 ? io_in_bits[111:104] : _GEN_1855; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2000 = 8'h7f == _T_28 ? io_in_bits[111:104] : _GEN_1856; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2001 = 8'h80 == _T_28 ? io_in_bits[111:104] : _GEN_1857; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2002 = 8'h81 == _T_28 ? io_in_bits[111:104] : _GEN_1858; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2003 = 8'h82 == _T_28 ? io_in_bits[111:104] : _GEN_1859; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2004 = 8'h83 == _T_28 ? io_in_bits[111:104] : _GEN_1860; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2005 = 8'h84 == _T_28 ? io_in_bits[111:104] : _GEN_1861; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2006 = 8'h85 == _T_28 ? io_in_bits[111:104] : _GEN_1862; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2007 = 8'h86 == _T_28 ? io_in_bits[111:104] : _GEN_1863; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2008 = 8'h87 == _T_28 ? io_in_bits[111:104] : _GEN_1864; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2009 = 8'h88 == _T_28 ? io_in_bits[111:104] : _GEN_1865; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2010 = 8'h89 == _T_28 ? io_in_bits[111:104] : _GEN_1866; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2011 = 8'h8a == _T_28 ? io_in_bits[111:104] : _GEN_1867; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2012 = 8'h8b == _T_28 ? io_in_bits[111:104] : _GEN_1868; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2013 = 8'h8c == _T_28 ? io_in_bits[111:104] : _GEN_1869; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2014 = 8'h8d == _T_28 ? io_in_bits[111:104] : _GEN_1870; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2015 = 8'h8e == _T_28 ? io_in_bits[111:104] : _GEN_1871; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _GEN_2016 = 8'h8f == _T_28 ? io_in_bits[111:104] : _GEN_1872; // @[WidthConverter.scala 67:{27,27}]
  wire [7:0] _T_30 = enqPtr + 8'he; // @[WidthConverter.scala 67:20]
  wire [7:0] _T_32 = enqPtr + 8'hf; // @[WidthConverter.scala 67:20]
  wire [7:0] _enqPtr_T_1 = enqPtr + 8'h10; // @[WidthConverter.scala 89:17]
  wire [7:0] _enqPtr_T_2 = _enqPtr_T_1 % 8'h90; // @[WidthConverter.scala 89:27]
  wire [7:0] _deqPtr_T_1 = deqPtr + 8'h9; // @[WidthConverter.scala 89:17]
  wire [7:0] _deqPtr_T_2 = _deqPtr_T_1 % 8'h90; // @[WidthConverter.scala 89:27]
  wire [7:0] _io_out_bits_T_3 = deqPtr + 8'h1; // @[WidthConverter.scala 84:26]
  wire [7:0] _io_out_bits_T_5 = deqPtr + 8'h2; // @[WidthConverter.scala 84:26]
  wire [7:0] _io_out_bits_T_7 = deqPtr + 8'h3; // @[WidthConverter.scala 84:26]
  wire [7:0] _io_out_bits_T_9 = deqPtr + 8'h4; // @[WidthConverter.scala 84:26]
  wire [7:0] _io_out_bits_T_11 = deqPtr + 8'h5; // @[WidthConverter.scala 84:26]
  wire [7:0] _io_out_bits_T_13 = deqPtr + 8'h6; // @[WidthConverter.scala 84:26]
  wire [7:0] _io_out_bits_T_15 = deqPtr + 8'h7; // @[WidthConverter.scala 84:26]
  wire [7:0] _io_out_bits_T_17 = deqPtr + 8'h8; // @[WidthConverter.scala 84:26]
  wire [7:0] _GEN_2452 = 8'h1 == _io_out_bits_T_3 ? arr_1 : arr_0; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2453 = 8'h2 == _io_out_bits_T_3 ? arr_2 : _GEN_2452; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2454 = 8'h3 == _io_out_bits_T_3 ? arr_3 : _GEN_2453; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2455 = 8'h4 == _io_out_bits_T_3 ? arr_4 : _GEN_2454; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2456 = 8'h5 == _io_out_bits_T_3 ? arr_5 : _GEN_2455; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2457 = 8'h6 == _io_out_bits_T_3 ? arr_6 : _GEN_2456; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2458 = 8'h7 == _io_out_bits_T_3 ? arr_7 : _GEN_2457; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2459 = 8'h8 == _io_out_bits_T_3 ? arr_8 : _GEN_2458; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2460 = 8'h9 == _io_out_bits_T_3 ? arr_9 : _GEN_2459; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2461 = 8'ha == _io_out_bits_T_3 ? arr_10 : _GEN_2460; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2462 = 8'hb == _io_out_bits_T_3 ? arr_11 : _GEN_2461; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2463 = 8'hc == _io_out_bits_T_3 ? arr_12 : _GEN_2462; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2464 = 8'hd == _io_out_bits_T_3 ? arr_13 : _GEN_2463; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2465 = 8'he == _io_out_bits_T_3 ? arr_14 : _GEN_2464; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2466 = 8'hf == _io_out_bits_T_3 ? arr_15 : _GEN_2465; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2467 = 8'h10 == _io_out_bits_T_3 ? arr_16 : _GEN_2466; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2468 = 8'h11 == _io_out_bits_T_3 ? arr_17 : _GEN_2467; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2469 = 8'h12 == _io_out_bits_T_3 ? arr_18 : _GEN_2468; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2470 = 8'h13 == _io_out_bits_T_3 ? arr_19 : _GEN_2469; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2471 = 8'h14 == _io_out_bits_T_3 ? arr_20 : _GEN_2470; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2472 = 8'h15 == _io_out_bits_T_3 ? arr_21 : _GEN_2471; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2473 = 8'h16 == _io_out_bits_T_3 ? arr_22 : _GEN_2472; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2474 = 8'h17 == _io_out_bits_T_3 ? arr_23 : _GEN_2473; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2475 = 8'h18 == _io_out_bits_T_3 ? arr_24 : _GEN_2474; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2476 = 8'h19 == _io_out_bits_T_3 ? arr_25 : _GEN_2475; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2477 = 8'h1a == _io_out_bits_T_3 ? arr_26 : _GEN_2476; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2478 = 8'h1b == _io_out_bits_T_3 ? arr_27 : _GEN_2477; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2479 = 8'h1c == _io_out_bits_T_3 ? arr_28 : _GEN_2478; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2480 = 8'h1d == _io_out_bits_T_3 ? arr_29 : _GEN_2479; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2481 = 8'h1e == _io_out_bits_T_3 ? arr_30 : _GEN_2480; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2482 = 8'h1f == _io_out_bits_T_3 ? arr_31 : _GEN_2481; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2483 = 8'h20 == _io_out_bits_T_3 ? arr_32 : _GEN_2482; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2484 = 8'h21 == _io_out_bits_T_3 ? arr_33 : _GEN_2483; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2485 = 8'h22 == _io_out_bits_T_3 ? arr_34 : _GEN_2484; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2486 = 8'h23 == _io_out_bits_T_3 ? arr_35 : _GEN_2485; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2487 = 8'h24 == _io_out_bits_T_3 ? arr_36 : _GEN_2486; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2488 = 8'h25 == _io_out_bits_T_3 ? arr_37 : _GEN_2487; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2489 = 8'h26 == _io_out_bits_T_3 ? arr_38 : _GEN_2488; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2490 = 8'h27 == _io_out_bits_T_3 ? arr_39 : _GEN_2489; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2491 = 8'h28 == _io_out_bits_T_3 ? arr_40 : _GEN_2490; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2492 = 8'h29 == _io_out_bits_T_3 ? arr_41 : _GEN_2491; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2493 = 8'h2a == _io_out_bits_T_3 ? arr_42 : _GEN_2492; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2494 = 8'h2b == _io_out_bits_T_3 ? arr_43 : _GEN_2493; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2495 = 8'h2c == _io_out_bits_T_3 ? arr_44 : _GEN_2494; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2496 = 8'h2d == _io_out_bits_T_3 ? arr_45 : _GEN_2495; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2497 = 8'h2e == _io_out_bits_T_3 ? arr_46 : _GEN_2496; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2498 = 8'h2f == _io_out_bits_T_3 ? arr_47 : _GEN_2497; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2499 = 8'h30 == _io_out_bits_T_3 ? arr_48 : _GEN_2498; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2500 = 8'h31 == _io_out_bits_T_3 ? arr_49 : _GEN_2499; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2501 = 8'h32 == _io_out_bits_T_3 ? arr_50 : _GEN_2500; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2502 = 8'h33 == _io_out_bits_T_3 ? arr_51 : _GEN_2501; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2503 = 8'h34 == _io_out_bits_T_3 ? arr_52 : _GEN_2502; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2504 = 8'h35 == _io_out_bits_T_3 ? arr_53 : _GEN_2503; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2505 = 8'h36 == _io_out_bits_T_3 ? arr_54 : _GEN_2504; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2506 = 8'h37 == _io_out_bits_T_3 ? arr_55 : _GEN_2505; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2507 = 8'h38 == _io_out_bits_T_3 ? arr_56 : _GEN_2506; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2508 = 8'h39 == _io_out_bits_T_3 ? arr_57 : _GEN_2507; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2509 = 8'h3a == _io_out_bits_T_3 ? arr_58 : _GEN_2508; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2510 = 8'h3b == _io_out_bits_T_3 ? arr_59 : _GEN_2509; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2511 = 8'h3c == _io_out_bits_T_3 ? arr_60 : _GEN_2510; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2512 = 8'h3d == _io_out_bits_T_3 ? arr_61 : _GEN_2511; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2513 = 8'h3e == _io_out_bits_T_3 ? arr_62 : _GEN_2512; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2514 = 8'h3f == _io_out_bits_T_3 ? arr_63 : _GEN_2513; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2515 = 8'h40 == _io_out_bits_T_3 ? arr_64 : _GEN_2514; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2516 = 8'h41 == _io_out_bits_T_3 ? arr_65 : _GEN_2515; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2517 = 8'h42 == _io_out_bits_T_3 ? arr_66 : _GEN_2516; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2518 = 8'h43 == _io_out_bits_T_3 ? arr_67 : _GEN_2517; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2519 = 8'h44 == _io_out_bits_T_3 ? arr_68 : _GEN_2518; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2520 = 8'h45 == _io_out_bits_T_3 ? arr_69 : _GEN_2519; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2521 = 8'h46 == _io_out_bits_T_3 ? arr_70 : _GEN_2520; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2522 = 8'h47 == _io_out_bits_T_3 ? arr_71 : _GEN_2521; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2523 = 8'h48 == _io_out_bits_T_3 ? arr_72 : _GEN_2522; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2524 = 8'h49 == _io_out_bits_T_3 ? arr_73 : _GEN_2523; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2525 = 8'h4a == _io_out_bits_T_3 ? arr_74 : _GEN_2524; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2526 = 8'h4b == _io_out_bits_T_3 ? arr_75 : _GEN_2525; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2527 = 8'h4c == _io_out_bits_T_3 ? arr_76 : _GEN_2526; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2528 = 8'h4d == _io_out_bits_T_3 ? arr_77 : _GEN_2527; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2529 = 8'h4e == _io_out_bits_T_3 ? arr_78 : _GEN_2528; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2530 = 8'h4f == _io_out_bits_T_3 ? arr_79 : _GEN_2529; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2531 = 8'h50 == _io_out_bits_T_3 ? arr_80 : _GEN_2530; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2532 = 8'h51 == _io_out_bits_T_3 ? arr_81 : _GEN_2531; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2533 = 8'h52 == _io_out_bits_T_3 ? arr_82 : _GEN_2532; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2534 = 8'h53 == _io_out_bits_T_3 ? arr_83 : _GEN_2533; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2535 = 8'h54 == _io_out_bits_T_3 ? arr_84 : _GEN_2534; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2536 = 8'h55 == _io_out_bits_T_3 ? arr_85 : _GEN_2535; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2537 = 8'h56 == _io_out_bits_T_3 ? arr_86 : _GEN_2536; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2538 = 8'h57 == _io_out_bits_T_3 ? arr_87 : _GEN_2537; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2539 = 8'h58 == _io_out_bits_T_3 ? arr_88 : _GEN_2538; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2540 = 8'h59 == _io_out_bits_T_3 ? arr_89 : _GEN_2539; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2541 = 8'h5a == _io_out_bits_T_3 ? arr_90 : _GEN_2540; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2542 = 8'h5b == _io_out_bits_T_3 ? arr_91 : _GEN_2541; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2543 = 8'h5c == _io_out_bits_T_3 ? arr_92 : _GEN_2542; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2544 = 8'h5d == _io_out_bits_T_3 ? arr_93 : _GEN_2543; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2545 = 8'h5e == _io_out_bits_T_3 ? arr_94 : _GEN_2544; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2546 = 8'h5f == _io_out_bits_T_3 ? arr_95 : _GEN_2545; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2547 = 8'h60 == _io_out_bits_T_3 ? arr_96 : _GEN_2546; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2548 = 8'h61 == _io_out_bits_T_3 ? arr_97 : _GEN_2547; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2549 = 8'h62 == _io_out_bits_T_3 ? arr_98 : _GEN_2548; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2550 = 8'h63 == _io_out_bits_T_3 ? arr_99 : _GEN_2549; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2551 = 8'h64 == _io_out_bits_T_3 ? arr_100 : _GEN_2550; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2552 = 8'h65 == _io_out_bits_T_3 ? arr_101 : _GEN_2551; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2553 = 8'h66 == _io_out_bits_T_3 ? arr_102 : _GEN_2552; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2554 = 8'h67 == _io_out_bits_T_3 ? arr_103 : _GEN_2553; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2555 = 8'h68 == _io_out_bits_T_3 ? arr_104 : _GEN_2554; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2556 = 8'h69 == _io_out_bits_T_3 ? arr_105 : _GEN_2555; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2557 = 8'h6a == _io_out_bits_T_3 ? arr_106 : _GEN_2556; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2558 = 8'h6b == _io_out_bits_T_3 ? arr_107 : _GEN_2557; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2559 = 8'h6c == _io_out_bits_T_3 ? arr_108 : _GEN_2558; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2560 = 8'h6d == _io_out_bits_T_3 ? arr_109 : _GEN_2559; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2561 = 8'h6e == _io_out_bits_T_3 ? arr_110 : _GEN_2560; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2562 = 8'h6f == _io_out_bits_T_3 ? arr_111 : _GEN_2561; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2563 = 8'h70 == _io_out_bits_T_3 ? arr_112 : _GEN_2562; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2564 = 8'h71 == _io_out_bits_T_3 ? arr_113 : _GEN_2563; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2565 = 8'h72 == _io_out_bits_T_3 ? arr_114 : _GEN_2564; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2566 = 8'h73 == _io_out_bits_T_3 ? arr_115 : _GEN_2565; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2567 = 8'h74 == _io_out_bits_T_3 ? arr_116 : _GEN_2566; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2568 = 8'h75 == _io_out_bits_T_3 ? arr_117 : _GEN_2567; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2569 = 8'h76 == _io_out_bits_T_3 ? arr_118 : _GEN_2568; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2570 = 8'h77 == _io_out_bits_T_3 ? arr_119 : _GEN_2569; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2571 = 8'h78 == _io_out_bits_T_3 ? arr_120 : _GEN_2570; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2572 = 8'h79 == _io_out_bits_T_3 ? arr_121 : _GEN_2571; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2573 = 8'h7a == _io_out_bits_T_3 ? arr_122 : _GEN_2572; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2574 = 8'h7b == _io_out_bits_T_3 ? arr_123 : _GEN_2573; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2575 = 8'h7c == _io_out_bits_T_3 ? arr_124 : _GEN_2574; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2576 = 8'h7d == _io_out_bits_T_3 ? arr_125 : _GEN_2575; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2577 = 8'h7e == _io_out_bits_T_3 ? arr_126 : _GEN_2576; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2578 = 8'h7f == _io_out_bits_T_3 ? arr_127 : _GEN_2577; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2579 = 8'h80 == _io_out_bits_T_3 ? arr_128 : _GEN_2578; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2580 = 8'h81 == _io_out_bits_T_3 ? arr_129 : _GEN_2579; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2581 = 8'h82 == _io_out_bits_T_3 ? arr_130 : _GEN_2580; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2582 = 8'h83 == _io_out_bits_T_3 ? arr_131 : _GEN_2581; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2583 = 8'h84 == _io_out_bits_T_3 ? arr_132 : _GEN_2582; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2584 = 8'h85 == _io_out_bits_T_3 ? arr_133 : _GEN_2583; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2585 = 8'h86 == _io_out_bits_T_3 ? arr_134 : _GEN_2584; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2586 = 8'h87 == _io_out_bits_T_3 ? arr_135 : _GEN_2585; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2587 = 8'h88 == _io_out_bits_T_3 ? arr_136 : _GEN_2586; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2588 = 8'h89 == _io_out_bits_T_3 ? arr_137 : _GEN_2587; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2589 = 8'h8a == _io_out_bits_T_3 ? arr_138 : _GEN_2588; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2590 = 8'h8b == _io_out_bits_T_3 ? arr_139 : _GEN_2589; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2591 = 8'h8c == _io_out_bits_T_3 ? arr_140 : _GEN_2590; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2592 = 8'h8d == _io_out_bits_T_3 ? arr_141 : _GEN_2591; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2593 = 8'h8e == _io_out_bits_T_3 ? arr_142 : _GEN_2592; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2594 = 8'h8f == _io_out_bits_T_3 ? arr_143 : _GEN_2593; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2596 = 8'h1 == _GEN_3747[7:0] ? arr_1 : arr_0; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2597 = 8'h2 == _GEN_3747[7:0] ? arr_2 : _GEN_2596; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2598 = 8'h3 == _GEN_3747[7:0] ? arr_3 : _GEN_2597; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2599 = 8'h4 == _GEN_3747[7:0] ? arr_4 : _GEN_2598; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2600 = 8'h5 == _GEN_3747[7:0] ? arr_5 : _GEN_2599; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2601 = 8'h6 == _GEN_3747[7:0] ? arr_6 : _GEN_2600; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2602 = 8'h7 == _GEN_3747[7:0] ? arr_7 : _GEN_2601; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2603 = 8'h8 == _GEN_3747[7:0] ? arr_8 : _GEN_2602; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2604 = 8'h9 == _GEN_3747[7:0] ? arr_9 : _GEN_2603; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2605 = 8'ha == _GEN_3747[7:0] ? arr_10 : _GEN_2604; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2606 = 8'hb == _GEN_3747[7:0] ? arr_11 : _GEN_2605; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2607 = 8'hc == _GEN_3747[7:0] ? arr_12 : _GEN_2606; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2608 = 8'hd == _GEN_3747[7:0] ? arr_13 : _GEN_2607; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2609 = 8'he == _GEN_3747[7:0] ? arr_14 : _GEN_2608; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2610 = 8'hf == _GEN_3747[7:0] ? arr_15 : _GEN_2609; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2611 = 8'h10 == _GEN_3747[7:0] ? arr_16 : _GEN_2610; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2612 = 8'h11 == _GEN_3747[7:0] ? arr_17 : _GEN_2611; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2613 = 8'h12 == _GEN_3747[7:0] ? arr_18 : _GEN_2612; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2614 = 8'h13 == _GEN_3747[7:0] ? arr_19 : _GEN_2613; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2615 = 8'h14 == _GEN_3747[7:0] ? arr_20 : _GEN_2614; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2616 = 8'h15 == _GEN_3747[7:0] ? arr_21 : _GEN_2615; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2617 = 8'h16 == _GEN_3747[7:0] ? arr_22 : _GEN_2616; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2618 = 8'h17 == _GEN_3747[7:0] ? arr_23 : _GEN_2617; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2619 = 8'h18 == _GEN_3747[7:0] ? arr_24 : _GEN_2618; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2620 = 8'h19 == _GEN_3747[7:0] ? arr_25 : _GEN_2619; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2621 = 8'h1a == _GEN_3747[7:0] ? arr_26 : _GEN_2620; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2622 = 8'h1b == _GEN_3747[7:0] ? arr_27 : _GEN_2621; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2623 = 8'h1c == _GEN_3747[7:0] ? arr_28 : _GEN_2622; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2624 = 8'h1d == _GEN_3747[7:0] ? arr_29 : _GEN_2623; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2625 = 8'h1e == _GEN_3747[7:0] ? arr_30 : _GEN_2624; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2626 = 8'h1f == _GEN_3747[7:0] ? arr_31 : _GEN_2625; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2627 = 8'h20 == _GEN_3747[7:0] ? arr_32 : _GEN_2626; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2628 = 8'h21 == _GEN_3747[7:0] ? arr_33 : _GEN_2627; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2629 = 8'h22 == _GEN_3747[7:0] ? arr_34 : _GEN_2628; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2630 = 8'h23 == _GEN_3747[7:0] ? arr_35 : _GEN_2629; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2631 = 8'h24 == _GEN_3747[7:0] ? arr_36 : _GEN_2630; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2632 = 8'h25 == _GEN_3747[7:0] ? arr_37 : _GEN_2631; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2633 = 8'h26 == _GEN_3747[7:0] ? arr_38 : _GEN_2632; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2634 = 8'h27 == _GEN_3747[7:0] ? arr_39 : _GEN_2633; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2635 = 8'h28 == _GEN_3747[7:0] ? arr_40 : _GEN_2634; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2636 = 8'h29 == _GEN_3747[7:0] ? arr_41 : _GEN_2635; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2637 = 8'h2a == _GEN_3747[7:0] ? arr_42 : _GEN_2636; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2638 = 8'h2b == _GEN_3747[7:0] ? arr_43 : _GEN_2637; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2639 = 8'h2c == _GEN_3747[7:0] ? arr_44 : _GEN_2638; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2640 = 8'h2d == _GEN_3747[7:0] ? arr_45 : _GEN_2639; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2641 = 8'h2e == _GEN_3747[7:0] ? arr_46 : _GEN_2640; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2642 = 8'h2f == _GEN_3747[7:0] ? arr_47 : _GEN_2641; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2643 = 8'h30 == _GEN_3747[7:0] ? arr_48 : _GEN_2642; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2644 = 8'h31 == _GEN_3747[7:0] ? arr_49 : _GEN_2643; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2645 = 8'h32 == _GEN_3747[7:0] ? arr_50 : _GEN_2644; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2646 = 8'h33 == _GEN_3747[7:0] ? arr_51 : _GEN_2645; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2647 = 8'h34 == _GEN_3747[7:0] ? arr_52 : _GEN_2646; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2648 = 8'h35 == _GEN_3747[7:0] ? arr_53 : _GEN_2647; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2649 = 8'h36 == _GEN_3747[7:0] ? arr_54 : _GEN_2648; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2650 = 8'h37 == _GEN_3747[7:0] ? arr_55 : _GEN_2649; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2651 = 8'h38 == _GEN_3747[7:0] ? arr_56 : _GEN_2650; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2652 = 8'h39 == _GEN_3747[7:0] ? arr_57 : _GEN_2651; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2653 = 8'h3a == _GEN_3747[7:0] ? arr_58 : _GEN_2652; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2654 = 8'h3b == _GEN_3747[7:0] ? arr_59 : _GEN_2653; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2655 = 8'h3c == _GEN_3747[7:0] ? arr_60 : _GEN_2654; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2656 = 8'h3d == _GEN_3747[7:0] ? arr_61 : _GEN_2655; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2657 = 8'h3e == _GEN_3747[7:0] ? arr_62 : _GEN_2656; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2658 = 8'h3f == _GEN_3747[7:0] ? arr_63 : _GEN_2657; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2659 = 8'h40 == _GEN_3747[7:0] ? arr_64 : _GEN_2658; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2660 = 8'h41 == _GEN_3747[7:0] ? arr_65 : _GEN_2659; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2661 = 8'h42 == _GEN_3747[7:0] ? arr_66 : _GEN_2660; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2662 = 8'h43 == _GEN_3747[7:0] ? arr_67 : _GEN_2661; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2663 = 8'h44 == _GEN_3747[7:0] ? arr_68 : _GEN_2662; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2664 = 8'h45 == _GEN_3747[7:0] ? arr_69 : _GEN_2663; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2665 = 8'h46 == _GEN_3747[7:0] ? arr_70 : _GEN_2664; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2666 = 8'h47 == _GEN_3747[7:0] ? arr_71 : _GEN_2665; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2667 = 8'h48 == _GEN_3747[7:0] ? arr_72 : _GEN_2666; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2668 = 8'h49 == _GEN_3747[7:0] ? arr_73 : _GEN_2667; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2669 = 8'h4a == _GEN_3747[7:0] ? arr_74 : _GEN_2668; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2670 = 8'h4b == _GEN_3747[7:0] ? arr_75 : _GEN_2669; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2671 = 8'h4c == _GEN_3747[7:0] ? arr_76 : _GEN_2670; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2672 = 8'h4d == _GEN_3747[7:0] ? arr_77 : _GEN_2671; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2673 = 8'h4e == _GEN_3747[7:0] ? arr_78 : _GEN_2672; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2674 = 8'h4f == _GEN_3747[7:0] ? arr_79 : _GEN_2673; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2675 = 8'h50 == _GEN_3747[7:0] ? arr_80 : _GEN_2674; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2676 = 8'h51 == _GEN_3747[7:0] ? arr_81 : _GEN_2675; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2677 = 8'h52 == _GEN_3747[7:0] ? arr_82 : _GEN_2676; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2678 = 8'h53 == _GEN_3747[7:0] ? arr_83 : _GEN_2677; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2679 = 8'h54 == _GEN_3747[7:0] ? arr_84 : _GEN_2678; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2680 = 8'h55 == _GEN_3747[7:0] ? arr_85 : _GEN_2679; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2681 = 8'h56 == _GEN_3747[7:0] ? arr_86 : _GEN_2680; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2682 = 8'h57 == _GEN_3747[7:0] ? arr_87 : _GEN_2681; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2683 = 8'h58 == _GEN_3747[7:0] ? arr_88 : _GEN_2682; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2684 = 8'h59 == _GEN_3747[7:0] ? arr_89 : _GEN_2683; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2685 = 8'h5a == _GEN_3747[7:0] ? arr_90 : _GEN_2684; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2686 = 8'h5b == _GEN_3747[7:0] ? arr_91 : _GEN_2685; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2687 = 8'h5c == _GEN_3747[7:0] ? arr_92 : _GEN_2686; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2688 = 8'h5d == _GEN_3747[7:0] ? arr_93 : _GEN_2687; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2689 = 8'h5e == _GEN_3747[7:0] ? arr_94 : _GEN_2688; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2690 = 8'h5f == _GEN_3747[7:0] ? arr_95 : _GEN_2689; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2691 = 8'h60 == _GEN_3747[7:0] ? arr_96 : _GEN_2690; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2692 = 8'h61 == _GEN_3747[7:0] ? arr_97 : _GEN_2691; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2693 = 8'h62 == _GEN_3747[7:0] ? arr_98 : _GEN_2692; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2694 = 8'h63 == _GEN_3747[7:0] ? arr_99 : _GEN_2693; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2695 = 8'h64 == _GEN_3747[7:0] ? arr_100 : _GEN_2694; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2696 = 8'h65 == _GEN_3747[7:0] ? arr_101 : _GEN_2695; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2697 = 8'h66 == _GEN_3747[7:0] ? arr_102 : _GEN_2696; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2698 = 8'h67 == _GEN_3747[7:0] ? arr_103 : _GEN_2697; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2699 = 8'h68 == _GEN_3747[7:0] ? arr_104 : _GEN_2698; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2700 = 8'h69 == _GEN_3747[7:0] ? arr_105 : _GEN_2699; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2701 = 8'h6a == _GEN_3747[7:0] ? arr_106 : _GEN_2700; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2702 = 8'h6b == _GEN_3747[7:0] ? arr_107 : _GEN_2701; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2703 = 8'h6c == _GEN_3747[7:0] ? arr_108 : _GEN_2702; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2704 = 8'h6d == _GEN_3747[7:0] ? arr_109 : _GEN_2703; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2705 = 8'h6e == _GEN_3747[7:0] ? arr_110 : _GEN_2704; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2706 = 8'h6f == _GEN_3747[7:0] ? arr_111 : _GEN_2705; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2707 = 8'h70 == _GEN_3747[7:0] ? arr_112 : _GEN_2706; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2708 = 8'h71 == _GEN_3747[7:0] ? arr_113 : _GEN_2707; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2709 = 8'h72 == _GEN_3747[7:0] ? arr_114 : _GEN_2708; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2710 = 8'h73 == _GEN_3747[7:0] ? arr_115 : _GEN_2709; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2711 = 8'h74 == _GEN_3747[7:0] ? arr_116 : _GEN_2710; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2712 = 8'h75 == _GEN_3747[7:0] ? arr_117 : _GEN_2711; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2713 = 8'h76 == _GEN_3747[7:0] ? arr_118 : _GEN_2712; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2714 = 8'h77 == _GEN_3747[7:0] ? arr_119 : _GEN_2713; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2715 = 8'h78 == _GEN_3747[7:0] ? arr_120 : _GEN_2714; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2716 = 8'h79 == _GEN_3747[7:0] ? arr_121 : _GEN_2715; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2717 = 8'h7a == _GEN_3747[7:0] ? arr_122 : _GEN_2716; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2718 = 8'h7b == _GEN_3747[7:0] ? arr_123 : _GEN_2717; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2719 = 8'h7c == _GEN_3747[7:0] ? arr_124 : _GEN_2718; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2720 = 8'h7d == _GEN_3747[7:0] ? arr_125 : _GEN_2719; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2721 = 8'h7e == _GEN_3747[7:0] ? arr_126 : _GEN_2720; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2722 = 8'h7f == _GEN_3747[7:0] ? arr_127 : _GEN_2721; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2723 = 8'h80 == _GEN_3747[7:0] ? arr_128 : _GEN_2722; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2724 = 8'h81 == _GEN_3747[7:0] ? arr_129 : _GEN_2723; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2725 = 8'h82 == _GEN_3747[7:0] ? arr_130 : _GEN_2724; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2726 = 8'h83 == _GEN_3747[7:0] ? arr_131 : _GEN_2725; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2727 = 8'h84 == _GEN_3747[7:0] ? arr_132 : _GEN_2726; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2728 = 8'h85 == _GEN_3747[7:0] ? arr_133 : _GEN_2727; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2729 = 8'h86 == _GEN_3747[7:0] ? arr_134 : _GEN_2728; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2730 = 8'h87 == _GEN_3747[7:0] ? arr_135 : _GEN_2729; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2731 = 8'h88 == _GEN_3747[7:0] ? arr_136 : _GEN_2730; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2732 = 8'h89 == _GEN_3747[7:0] ? arr_137 : _GEN_2731; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2733 = 8'h8a == _GEN_3747[7:0] ? arr_138 : _GEN_2732; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2734 = 8'h8b == _GEN_3747[7:0] ? arr_139 : _GEN_2733; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2735 = 8'h8c == _GEN_3747[7:0] ? arr_140 : _GEN_2734; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2736 = 8'h8d == _GEN_3747[7:0] ? arr_141 : _GEN_2735; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2737 = 8'h8e == _GEN_3747[7:0] ? arr_142 : _GEN_2736; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2738 = 8'h8f == _GEN_3747[7:0] ? arr_143 : _GEN_2737; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2740 = 8'h1 == _io_out_bits_T_7 ? arr_1 : arr_0; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2741 = 8'h2 == _io_out_bits_T_7 ? arr_2 : _GEN_2740; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2742 = 8'h3 == _io_out_bits_T_7 ? arr_3 : _GEN_2741; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2743 = 8'h4 == _io_out_bits_T_7 ? arr_4 : _GEN_2742; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2744 = 8'h5 == _io_out_bits_T_7 ? arr_5 : _GEN_2743; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2745 = 8'h6 == _io_out_bits_T_7 ? arr_6 : _GEN_2744; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2746 = 8'h7 == _io_out_bits_T_7 ? arr_7 : _GEN_2745; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2747 = 8'h8 == _io_out_bits_T_7 ? arr_8 : _GEN_2746; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2748 = 8'h9 == _io_out_bits_T_7 ? arr_9 : _GEN_2747; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2749 = 8'ha == _io_out_bits_T_7 ? arr_10 : _GEN_2748; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2750 = 8'hb == _io_out_bits_T_7 ? arr_11 : _GEN_2749; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2751 = 8'hc == _io_out_bits_T_7 ? arr_12 : _GEN_2750; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2752 = 8'hd == _io_out_bits_T_7 ? arr_13 : _GEN_2751; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2753 = 8'he == _io_out_bits_T_7 ? arr_14 : _GEN_2752; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2754 = 8'hf == _io_out_bits_T_7 ? arr_15 : _GEN_2753; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2755 = 8'h10 == _io_out_bits_T_7 ? arr_16 : _GEN_2754; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2756 = 8'h11 == _io_out_bits_T_7 ? arr_17 : _GEN_2755; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2757 = 8'h12 == _io_out_bits_T_7 ? arr_18 : _GEN_2756; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2758 = 8'h13 == _io_out_bits_T_7 ? arr_19 : _GEN_2757; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2759 = 8'h14 == _io_out_bits_T_7 ? arr_20 : _GEN_2758; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2760 = 8'h15 == _io_out_bits_T_7 ? arr_21 : _GEN_2759; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2761 = 8'h16 == _io_out_bits_T_7 ? arr_22 : _GEN_2760; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2762 = 8'h17 == _io_out_bits_T_7 ? arr_23 : _GEN_2761; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2763 = 8'h18 == _io_out_bits_T_7 ? arr_24 : _GEN_2762; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2764 = 8'h19 == _io_out_bits_T_7 ? arr_25 : _GEN_2763; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2765 = 8'h1a == _io_out_bits_T_7 ? arr_26 : _GEN_2764; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2766 = 8'h1b == _io_out_bits_T_7 ? arr_27 : _GEN_2765; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2767 = 8'h1c == _io_out_bits_T_7 ? arr_28 : _GEN_2766; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2768 = 8'h1d == _io_out_bits_T_7 ? arr_29 : _GEN_2767; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2769 = 8'h1e == _io_out_bits_T_7 ? arr_30 : _GEN_2768; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2770 = 8'h1f == _io_out_bits_T_7 ? arr_31 : _GEN_2769; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2771 = 8'h20 == _io_out_bits_T_7 ? arr_32 : _GEN_2770; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2772 = 8'h21 == _io_out_bits_T_7 ? arr_33 : _GEN_2771; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2773 = 8'h22 == _io_out_bits_T_7 ? arr_34 : _GEN_2772; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2774 = 8'h23 == _io_out_bits_T_7 ? arr_35 : _GEN_2773; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2775 = 8'h24 == _io_out_bits_T_7 ? arr_36 : _GEN_2774; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2776 = 8'h25 == _io_out_bits_T_7 ? arr_37 : _GEN_2775; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2777 = 8'h26 == _io_out_bits_T_7 ? arr_38 : _GEN_2776; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2778 = 8'h27 == _io_out_bits_T_7 ? arr_39 : _GEN_2777; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2779 = 8'h28 == _io_out_bits_T_7 ? arr_40 : _GEN_2778; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2780 = 8'h29 == _io_out_bits_T_7 ? arr_41 : _GEN_2779; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2781 = 8'h2a == _io_out_bits_T_7 ? arr_42 : _GEN_2780; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2782 = 8'h2b == _io_out_bits_T_7 ? arr_43 : _GEN_2781; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2783 = 8'h2c == _io_out_bits_T_7 ? arr_44 : _GEN_2782; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2784 = 8'h2d == _io_out_bits_T_7 ? arr_45 : _GEN_2783; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2785 = 8'h2e == _io_out_bits_T_7 ? arr_46 : _GEN_2784; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2786 = 8'h2f == _io_out_bits_T_7 ? arr_47 : _GEN_2785; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2787 = 8'h30 == _io_out_bits_T_7 ? arr_48 : _GEN_2786; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2788 = 8'h31 == _io_out_bits_T_7 ? arr_49 : _GEN_2787; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2789 = 8'h32 == _io_out_bits_T_7 ? arr_50 : _GEN_2788; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2790 = 8'h33 == _io_out_bits_T_7 ? arr_51 : _GEN_2789; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2791 = 8'h34 == _io_out_bits_T_7 ? arr_52 : _GEN_2790; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2792 = 8'h35 == _io_out_bits_T_7 ? arr_53 : _GEN_2791; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2793 = 8'h36 == _io_out_bits_T_7 ? arr_54 : _GEN_2792; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2794 = 8'h37 == _io_out_bits_T_7 ? arr_55 : _GEN_2793; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2795 = 8'h38 == _io_out_bits_T_7 ? arr_56 : _GEN_2794; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2796 = 8'h39 == _io_out_bits_T_7 ? arr_57 : _GEN_2795; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2797 = 8'h3a == _io_out_bits_T_7 ? arr_58 : _GEN_2796; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2798 = 8'h3b == _io_out_bits_T_7 ? arr_59 : _GEN_2797; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2799 = 8'h3c == _io_out_bits_T_7 ? arr_60 : _GEN_2798; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2800 = 8'h3d == _io_out_bits_T_7 ? arr_61 : _GEN_2799; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2801 = 8'h3e == _io_out_bits_T_7 ? arr_62 : _GEN_2800; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2802 = 8'h3f == _io_out_bits_T_7 ? arr_63 : _GEN_2801; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2803 = 8'h40 == _io_out_bits_T_7 ? arr_64 : _GEN_2802; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2804 = 8'h41 == _io_out_bits_T_7 ? arr_65 : _GEN_2803; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2805 = 8'h42 == _io_out_bits_T_7 ? arr_66 : _GEN_2804; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2806 = 8'h43 == _io_out_bits_T_7 ? arr_67 : _GEN_2805; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2807 = 8'h44 == _io_out_bits_T_7 ? arr_68 : _GEN_2806; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2808 = 8'h45 == _io_out_bits_T_7 ? arr_69 : _GEN_2807; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2809 = 8'h46 == _io_out_bits_T_7 ? arr_70 : _GEN_2808; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2810 = 8'h47 == _io_out_bits_T_7 ? arr_71 : _GEN_2809; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2811 = 8'h48 == _io_out_bits_T_7 ? arr_72 : _GEN_2810; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2812 = 8'h49 == _io_out_bits_T_7 ? arr_73 : _GEN_2811; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2813 = 8'h4a == _io_out_bits_T_7 ? arr_74 : _GEN_2812; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2814 = 8'h4b == _io_out_bits_T_7 ? arr_75 : _GEN_2813; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2815 = 8'h4c == _io_out_bits_T_7 ? arr_76 : _GEN_2814; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2816 = 8'h4d == _io_out_bits_T_7 ? arr_77 : _GEN_2815; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2817 = 8'h4e == _io_out_bits_T_7 ? arr_78 : _GEN_2816; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2818 = 8'h4f == _io_out_bits_T_7 ? arr_79 : _GEN_2817; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2819 = 8'h50 == _io_out_bits_T_7 ? arr_80 : _GEN_2818; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2820 = 8'h51 == _io_out_bits_T_7 ? arr_81 : _GEN_2819; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2821 = 8'h52 == _io_out_bits_T_7 ? arr_82 : _GEN_2820; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2822 = 8'h53 == _io_out_bits_T_7 ? arr_83 : _GEN_2821; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2823 = 8'h54 == _io_out_bits_T_7 ? arr_84 : _GEN_2822; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2824 = 8'h55 == _io_out_bits_T_7 ? arr_85 : _GEN_2823; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2825 = 8'h56 == _io_out_bits_T_7 ? arr_86 : _GEN_2824; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2826 = 8'h57 == _io_out_bits_T_7 ? arr_87 : _GEN_2825; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2827 = 8'h58 == _io_out_bits_T_7 ? arr_88 : _GEN_2826; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2828 = 8'h59 == _io_out_bits_T_7 ? arr_89 : _GEN_2827; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2829 = 8'h5a == _io_out_bits_T_7 ? arr_90 : _GEN_2828; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2830 = 8'h5b == _io_out_bits_T_7 ? arr_91 : _GEN_2829; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2831 = 8'h5c == _io_out_bits_T_7 ? arr_92 : _GEN_2830; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2832 = 8'h5d == _io_out_bits_T_7 ? arr_93 : _GEN_2831; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2833 = 8'h5e == _io_out_bits_T_7 ? arr_94 : _GEN_2832; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2834 = 8'h5f == _io_out_bits_T_7 ? arr_95 : _GEN_2833; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2835 = 8'h60 == _io_out_bits_T_7 ? arr_96 : _GEN_2834; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2836 = 8'h61 == _io_out_bits_T_7 ? arr_97 : _GEN_2835; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2837 = 8'h62 == _io_out_bits_T_7 ? arr_98 : _GEN_2836; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2838 = 8'h63 == _io_out_bits_T_7 ? arr_99 : _GEN_2837; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2839 = 8'h64 == _io_out_bits_T_7 ? arr_100 : _GEN_2838; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2840 = 8'h65 == _io_out_bits_T_7 ? arr_101 : _GEN_2839; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2841 = 8'h66 == _io_out_bits_T_7 ? arr_102 : _GEN_2840; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2842 = 8'h67 == _io_out_bits_T_7 ? arr_103 : _GEN_2841; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2843 = 8'h68 == _io_out_bits_T_7 ? arr_104 : _GEN_2842; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2844 = 8'h69 == _io_out_bits_T_7 ? arr_105 : _GEN_2843; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2845 = 8'h6a == _io_out_bits_T_7 ? arr_106 : _GEN_2844; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2846 = 8'h6b == _io_out_bits_T_7 ? arr_107 : _GEN_2845; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2847 = 8'h6c == _io_out_bits_T_7 ? arr_108 : _GEN_2846; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2848 = 8'h6d == _io_out_bits_T_7 ? arr_109 : _GEN_2847; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2849 = 8'h6e == _io_out_bits_T_7 ? arr_110 : _GEN_2848; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2850 = 8'h6f == _io_out_bits_T_7 ? arr_111 : _GEN_2849; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2851 = 8'h70 == _io_out_bits_T_7 ? arr_112 : _GEN_2850; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2852 = 8'h71 == _io_out_bits_T_7 ? arr_113 : _GEN_2851; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2853 = 8'h72 == _io_out_bits_T_7 ? arr_114 : _GEN_2852; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2854 = 8'h73 == _io_out_bits_T_7 ? arr_115 : _GEN_2853; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2855 = 8'h74 == _io_out_bits_T_7 ? arr_116 : _GEN_2854; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2856 = 8'h75 == _io_out_bits_T_7 ? arr_117 : _GEN_2855; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2857 = 8'h76 == _io_out_bits_T_7 ? arr_118 : _GEN_2856; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2858 = 8'h77 == _io_out_bits_T_7 ? arr_119 : _GEN_2857; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2859 = 8'h78 == _io_out_bits_T_7 ? arr_120 : _GEN_2858; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2860 = 8'h79 == _io_out_bits_T_7 ? arr_121 : _GEN_2859; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2861 = 8'h7a == _io_out_bits_T_7 ? arr_122 : _GEN_2860; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2862 = 8'h7b == _io_out_bits_T_7 ? arr_123 : _GEN_2861; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2863 = 8'h7c == _io_out_bits_T_7 ? arr_124 : _GEN_2862; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2864 = 8'h7d == _io_out_bits_T_7 ? arr_125 : _GEN_2863; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2865 = 8'h7e == _io_out_bits_T_7 ? arr_126 : _GEN_2864; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2866 = 8'h7f == _io_out_bits_T_7 ? arr_127 : _GEN_2865; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2867 = 8'h80 == _io_out_bits_T_7 ? arr_128 : _GEN_2866; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2868 = 8'h81 == _io_out_bits_T_7 ? arr_129 : _GEN_2867; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2869 = 8'h82 == _io_out_bits_T_7 ? arr_130 : _GEN_2868; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2870 = 8'h83 == _io_out_bits_T_7 ? arr_131 : _GEN_2869; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2871 = 8'h84 == _io_out_bits_T_7 ? arr_132 : _GEN_2870; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2872 = 8'h85 == _io_out_bits_T_7 ? arr_133 : _GEN_2871; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2873 = 8'h86 == _io_out_bits_T_7 ? arr_134 : _GEN_2872; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2874 = 8'h87 == _io_out_bits_T_7 ? arr_135 : _GEN_2873; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2875 = 8'h88 == _io_out_bits_T_7 ? arr_136 : _GEN_2874; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2876 = 8'h89 == _io_out_bits_T_7 ? arr_137 : _GEN_2875; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2877 = 8'h8a == _io_out_bits_T_7 ? arr_138 : _GEN_2876; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2878 = 8'h8b == _io_out_bits_T_7 ? arr_139 : _GEN_2877; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2879 = 8'h8c == _io_out_bits_T_7 ? arr_140 : _GEN_2878; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2880 = 8'h8d == _io_out_bits_T_7 ? arr_141 : _GEN_2879; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2881 = 8'h8e == _io_out_bits_T_7 ? arr_142 : _GEN_2880; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2882 = 8'h8f == _io_out_bits_T_7 ? arr_143 : _GEN_2881; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2884 = 8'h1 == _io_out_bits_T_5 ? arr_1 : arr_0; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2885 = 8'h2 == _io_out_bits_T_5 ? arr_2 : _GEN_2884; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2886 = 8'h3 == _io_out_bits_T_5 ? arr_3 : _GEN_2885; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2887 = 8'h4 == _io_out_bits_T_5 ? arr_4 : _GEN_2886; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2888 = 8'h5 == _io_out_bits_T_5 ? arr_5 : _GEN_2887; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2889 = 8'h6 == _io_out_bits_T_5 ? arr_6 : _GEN_2888; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2890 = 8'h7 == _io_out_bits_T_5 ? arr_7 : _GEN_2889; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2891 = 8'h8 == _io_out_bits_T_5 ? arr_8 : _GEN_2890; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2892 = 8'h9 == _io_out_bits_T_5 ? arr_9 : _GEN_2891; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2893 = 8'ha == _io_out_bits_T_5 ? arr_10 : _GEN_2892; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2894 = 8'hb == _io_out_bits_T_5 ? arr_11 : _GEN_2893; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2895 = 8'hc == _io_out_bits_T_5 ? arr_12 : _GEN_2894; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2896 = 8'hd == _io_out_bits_T_5 ? arr_13 : _GEN_2895; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2897 = 8'he == _io_out_bits_T_5 ? arr_14 : _GEN_2896; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2898 = 8'hf == _io_out_bits_T_5 ? arr_15 : _GEN_2897; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2899 = 8'h10 == _io_out_bits_T_5 ? arr_16 : _GEN_2898; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2900 = 8'h11 == _io_out_bits_T_5 ? arr_17 : _GEN_2899; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2901 = 8'h12 == _io_out_bits_T_5 ? arr_18 : _GEN_2900; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2902 = 8'h13 == _io_out_bits_T_5 ? arr_19 : _GEN_2901; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2903 = 8'h14 == _io_out_bits_T_5 ? arr_20 : _GEN_2902; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2904 = 8'h15 == _io_out_bits_T_5 ? arr_21 : _GEN_2903; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2905 = 8'h16 == _io_out_bits_T_5 ? arr_22 : _GEN_2904; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2906 = 8'h17 == _io_out_bits_T_5 ? arr_23 : _GEN_2905; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2907 = 8'h18 == _io_out_bits_T_5 ? arr_24 : _GEN_2906; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2908 = 8'h19 == _io_out_bits_T_5 ? arr_25 : _GEN_2907; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2909 = 8'h1a == _io_out_bits_T_5 ? arr_26 : _GEN_2908; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2910 = 8'h1b == _io_out_bits_T_5 ? arr_27 : _GEN_2909; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2911 = 8'h1c == _io_out_bits_T_5 ? arr_28 : _GEN_2910; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2912 = 8'h1d == _io_out_bits_T_5 ? arr_29 : _GEN_2911; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2913 = 8'h1e == _io_out_bits_T_5 ? arr_30 : _GEN_2912; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2914 = 8'h1f == _io_out_bits_T_5 ? arr_31 : _GEN_2913; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2915 = 8'h20 == _io_out_bits_T_5 ? arr_32 : _GEN_2914; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2916 = 8'h21 == _io_out_bits_T_5 ? arr_33 : _GEN_2915; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2917 = 8'h22 == _io_out_bits_T_5 ? arr_34 : _GEN_2916; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2918 = 8'h23 == _io_out_bits_T_5 ? arr_35 : _GEN_2917; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2919 = 8'h24 == _io_out_bits_T_5 ? arr_36 : _GEN_2918; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2920 = 8'h25 == _io_out_bits_T_5 ? arr_37 : _GEN_2919; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2921 = 8'h26 == _io_out_bits_T_5 ? arr_38 : _GEN_2920; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2922 = 8'h27 == _io_out_bits_T_5 ? arr_39 : _GEN_2921; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2923 = 8'h28 == _io_out_bits_T_5 ? arr_40 : _GEN_2922; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2924 = 8'h29 == _io_out_bits_T_5 ? arr_41 : _GEN_2923; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2925 = 8'h2a == _io_out_bits_T_5 ? arr_42 : _GEN_2924; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2926 = 8'h2b == _io_out_bits_T_5 ? arr_43 : _GEN_2925; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2927 = 8'h2c == _io_out_bits_T_5 ? arr_44 : _GEN_2926; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2928 = 8'h2d == _io_out_bits_T_5 ? arr_45 : _GEN_2927; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2929 = 8'h2e == _io_out_bits_T_5 ? arr_46 : _GEN_2928; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2930 = 8'h2f == _io_out_bits_T_5 ? arr_47 : _GEN_2929; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2931 = 8'h30 == _io_out_bits_T_5 ? arr_48 : _GEN_2930; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2932 = 8'h31 == _io_out_bits_T_5 ? arr_49 : _GEN_2931; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2933 = 8'h32 == _io_out_bits_T_5 ? arr_50 : _GEN_2932; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2934 = 8'h33 == _io_out_bits_T_5 ? arr_51 : _GEN_2933; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2935 = 8'h34 == _io_out_bits_T_5 ? arr_52 : _GEN_2934; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2936 = 8'h35 == _io_out_bits_T_5 ? arr_53 : _GEN_2935; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2937 = 8'h36 == _io_out_bits_T_5 ? arr_54 : _GEN_2936; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2938 = 8'h37 == _io_out_bits_T_5 ? arr_55 : _GEN_2937; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2939 = 8'h38 == _io_out_bits_T_5 ? arr_56 : _GEN_2938; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2940 = 8'h39 == _io_out_bits_T_5 ? arr_57 : _GEN_2939; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2941 = 8'h3a == _io_out_bits_T_5 ? arr_58 : _GEN_2940; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2942 = 8'h3b == _io_out_bits_T_5 ? arr_59 : _GEN_2941; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2943 = 8'h3c == _io_out_bits_T_5 ? arr_60 : _GEN_2942; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2944 = 8'h3d == _io_out_bits_T_5 ? arr_61 : _GEN_2943; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2945 = 8'h3e == _io_out_bits_T_5 ? arr_62 : _GEN_2944; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2946 = 8'h3f == _io_out_bits_T_5 ? arr_63 : _GEN_2945; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2947 = 8'h40 == _io_out_bits_T_5 ? arr_64 : _GEN_2946; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2948 = 8'h41 == _io_out_bits_T_5 ? arr_65 : _GEN_2947; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2949 = 8'h42 == _io_out_bits_T_5 ? arr_66 : _GEN_2948; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2950 = 8'h43 == _io_out_bits_T_5 ? arr_67 : _GEN_2949; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2951 = 8'h44 == _io_out_bits_T_5 ? arr_68 : _GEN_2950; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2952 = 8'h45 == _io_out_bits_T_5 ? arr_69 : _GEN_2951; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2953 = 8'h46 == _io_out_bits_T_5 ? arr_70 : _GEN_2952; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2954 = 8'h47 == _io_out_bits_T_5 ? arr_71 : _GEN_2953; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2955 = 8'h48 == _io_out_bits_T_5 ? arr_72 : _GEN_2954; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2956 = 8'h49 == _io_out_bits_T_5 ? arr_73 : _GEN_2955; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2957 = 8'h4a == _io_out_bits_T_5 ? arr_74 : _GEN_2956; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2958 = 8'h4b == _io_out_bits_T_5 ? arr_75 : _GEN_2957; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2959 = 8'h4c == _io_out_bits_T_5 ? arr_76 : _GEN_2958; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2960 = 8'h4d == _io_out_bits_T_5 ? arr_77 : _GEN_2959; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2961 = 8'h4e == _io_out_bits_T_5 ? arr_78 : _GEN_2960; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2962 = 8'h4f == _io_out_bits_T_5 ? arr_79 : _GEN_2961; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2963 = 8'h50 == _io_out_bits_T_5 ? arr_80 : _GEN_2962; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2964 = 8'h51 == _io_out_bits_T_5 ? arr_81 : _GEN_2963; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2965 = 8'h52 == _io_out_bits_T_5 ? arr_82 : _GEN_2964; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2966 = 8'h53 == _io_out_bits_T_5 ? arr_83 : _GEN_2965; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2967 = 8'h54 == _io_out_bits_T_5 ? arr_84 : _GEN_2966; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2968 = 8'h55 == _io_out_bits_T_5 ? arr_85 : _GEN_2967; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2969 = 8'h56 == _io_out_bits_T_5 ? arr_86 : _GEN_2968; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2970 = 8'h57 == _io_out_bits_T_5 ? arr_87 : _GEN_2969; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2971 = 8'h58 == _io_out_bits_T_5 ? arr_88 : _GEN_2970; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2972 = 8'h59 == _io_out_bits_T_5 ? arr_89 : _GEN_2971; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2973 = 8'h5a == _io_out_bits_T_5 ? arr_90 : _GEN_2972; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2974 = 8'h5b == _io_out_bits_T_5 ? arr_91 : _GEN_2973; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2975 = 8'h5c == _io_out_bits_T_5 ? arr_92 : _GEN_2974; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2976 = 8'h5d == _io_out_bits_T_5 ? arr_93 : _GEN_2975; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2977 = 8'h5e == _io_out_bits_T_5 ? arr_94 : _GEN_2976; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2978 = 8'h5f == _io_out_bits_T_5 ? arr_95 : _GEN_2977; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2979 = 8'h60 == _io_out_bits_T_5 ? arr_96 : _GEN_2978; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2980 = 8'h61 == _io_out_bits_T_5 ? arr_97 : _GEN_2979; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2981 = 8'h62 == _io_out_bits_T_5 ? arr_98 : _GEN_2980; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2982 = 8'h63 == _io_out_bits_T_5 ? arr_99 : _GEN_2981; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2983 = 8'h64 == _io_out_bits_T_5 ? arr_100 : _GEN_2982; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2984 = 8'h65 == _io_out_bits_T_5 ? arr_101 : _GEN_2983; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2985 = 8'h66 == _io_out_bits_T_5 ? arr_102 : _GEN_2984; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2986 = 8'h67 == _io_out_bits_T_5 ? arr_103 : _GEN_2985; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2987 = 8'h68 == _io_out_bits_T_5 ? arr_104 : _GEN_2986; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2988 = 8'h69 == _io_out_bits_T_5 ? arr_105 : _GEN_2987; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2989 = 8'h6a == _io_out_bits_T_5 ? arr_106 : _GEN_2988; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2990 = 8'h6b == _io_out_bits_T_5 ? arr_107 : _GEN_2989; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2991 = 8'h6c == _io_out_bits_T_5 ? arr_108 : _GEN_2990; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2992 = 8'h6d == _io_out_bits_T_5 ? arr_109 : _GEN_2991; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2993 = 8'h6e == _io_out_bits_T_5 ? arr_110 : _GEN_2992; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2994 = 8'h6f == _io_out_bits_T_5 ? arr_111 : _GEN_2993; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2995 = 8'h70 == _io_out_bits_T_5 ? arr_112 : _GEN_2994; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2996 = 8'h71 == _io_out_bits_T_5 ? arr_113 : _GEN_2995; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2997 = 8'h72 == _io_out_bits_T_5 ? arr_114 : _GEN_2996; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2998 = 8'h73 == _io_out_bits_T_5 ? arr_115 : _GEN_2997; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_2999 = 8'h74 == _io_out_bits_T_5 ? arr_116 : _GEN_2998; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3000 = 8'h75 == _io_out_bits_T_5 ? arr_117 : _GEN_2999; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3001 = 8'h76 == _io_out_bits_T_5 ? arr_118 : _GEN_3000; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3002 = 8'h77 == _io_out_bits_T_5 ? arr_119 : _GEN_3001; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3003 = 8'h78 == _io_out_bits_T_5 ? arr_120 : _GEN_3002; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3004 = 8'h79 == _io_out_bits_T_5 ? arr_121 : _GEN_3003; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3005 = 8'h7a == _io_out_bits_T_5 ? arr_122 : _GEN_3004; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3006 = 8'h7b == _io_out_bits_T_5 ? arr_123 : _GEN_3005; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3007 = 8'h7c == _io_out_bits_T_5 ? arr_124 : _GEN_3006; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3008 = 8'h7d == _io_out_bits_T_5 ? arr_125 : _GEN_3007; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3009 = 8'h7e == _io_out_bits_T_5 ? arr_126 : _GEN_3008; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3010 = 8'h7f == _io_out_bits_T_5 ? arr_127 : _GEN_3009; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3011 = 8'h80 == _io_out_bits_T_5 ? arr_128 : _GEN_3010; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3012 = 8'h81 == _io_out_bits_T_5 ? arr_129 : _GEN_3011; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3013 = 8'h82 == _io_out_bits_T_5 ? arr_130 : _GEN_3012; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3014 = 8'h83 == _io_out_bits_T_5 ? arr_131 : _GEN_3013; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3015 = 8'h84 == _io_out_bits_T_5 ? arr_132 : _GEN_3014; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3016 = 8'h85 == _io_out_bits_T_5 ? arr_133 : _GEN_3015; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3017 = 8'h86 == _io_out_bits_T_5 ? arr_134 : _GEN_3016; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3018 = 8'h87 == _io_out_bits_T_5 ? arr_135 : _GEN_3017; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3019 = 8'h88 == _io_out_bits_T_5 ? arr_136 : _GEN_3018; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3020 = 8'h89 == _io_out_bits_T_5 ? arr_137 : _GEN_3019; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3021 = 8'h8a == _io_out_bits_T_5 ? arr_138 : _GEN_3020; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3022 = 8'h8b == _io_out_bits_T_5 ? arr_139 : _GEN_3021; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3023 = 8'h8c == _io_out_bits_T_5 ? arr_140 : _GEN_3022; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3024 = 8'h8d == _io_out_bits_T_5 ? arr_141 : _GEN_3023; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3025 = 8'h8e == _io_out_bits_T_5 ? arr_142 : _GEN_3024; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3026 = 8'h8f == _io_out_bits_T_5 ? arr_143 : _GEN_3025; // @[Cat.scala 31:{58,58}]
  wire [31:0] io_out_bits_lo = {_GEN_2882,_GEN_3026,_GEN_2594,_GEN_2738}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_3028 = 8'h1 == _io_out_bits_T_11 ? arr_1 : arr_0; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3029 = 8'h2 == _io_out_bits_T_11 ? arr_2 : _GEN_3028; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3030 = 8'h3 == _io_out_bits_T_11 ? arr_3 : _GEN_3029; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3031 = 8'h4 == _io_out_bits_T_11 ? arr_4 : _GEN_3030; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3032 = 8'h5 == _io_out_bits_T_11 ? arr_5 : _GEN_3031; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3033 = 8'h6 == _io_out_bits_T_11 ? arr_6 : _GEN_3032; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3034 = 8'h7 == _io_out_bits_T_11 ? arr_7 : _GEN_3033; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3035 = 8'h8 == _io_out_bits_T_11 ? arr_8 : _GEN_3034; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3036 = 8'h9 == _io_out_bits_T_11 ? arr_9 : _GEN_3035; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3037 = 8'ha == _io_out_bits_T_11 ? arr_10 : _GEN_3036; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3038 = 8'hb == _io_out_bits_T_11 ? arr_11 : _GEN_3037; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3039 = 8'hc == _io_out_bits_T_11 ? arr_12 : _GEN_3038; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3040 = 8'hd == _io_out_bits_T_11 ? arr_13 : _GEN_3039; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3041 = 8'he == _io_out_bits_T_11 ? arr_14 : _GEN_3040; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3042 = 8'hf == _io_out_bits_T_11 ? arr_15 : _GEN_3041; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3043 = 8'h10 == _io_out_bits_T_11 ? arr_16 : _GEN_3042; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3044 = 8'h11 == _io_out_bits_T_11 ? arr_17 : _GEN_3043; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3045 = 8'h12 == _io_out_bits_T_11 ? arr_18 : _GEN_3044; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3046 = 8'h13 == _io_out_bits_T_11 ? arr_19 : _GEN_3045; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3047 = 8'h14 == _io_out_bits_T_11 ? arr_20 : _GEN_3046; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3048 = 8'h15 == _io_out_bits_T_11 ? arr_21 : _GEN_3047; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3049 = 8'h16 == _io_out_bits_T_11 ? arr_22 : _GEN_3048; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3050 = 8'h17 == _io_out_bits_T_11 ? arr_23 : _GEN_3049; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3051 = 8'h18 == _io_out_bits_T_11 ? arr_24 : _GEN_3050; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3052 = 8'h19 == _io_out_bits_T_11 ? arr_25 : _GEN_3051; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3053 = 8'h1a == _io_out_bits_T_11 ? arr_26 : _GEN_3052; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3054 = 8'h1b == _io_out_bits_T_11 ? arr_27 : _GEN_3053; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3055 = 8'h1c == _io_out_bits_T_11 ? arr_28 : _GEN_3054; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3056 = 8'h1d == _io_out_bits_T_11 ? arr_29 : _GEN_3055; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3057 = 8'h1e == _io_out_bits_T_11 ? arr_30 : _GEN_3056; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3058 = 8'h1f == _io_out_bits_T_11 ? arr_31 : _GEN_3057; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3059 = 8'h20 == _io_out_bits_T_11 ? arr_32 : _GEN_3058; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3060 = 8'h21 == _io_out_bits_T_11 ? arr_33 : _GEN_3059; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3061 = 8'h22 == _io_out_bits_T_11 ? arr_34 : _GEN_3060; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3062 = 8'h23 == _io_out_bits_T_11 ? arr_35 : _GEN_3061; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3063 = 8'h24 == _io_out_bits_T_11 ? arr_36 : _GEN_3062; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3064 = 8'h25 == _io_out_bits_T_11 ? arr_37 : _GEN_3063; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3065 = 8'h26 == _io_out_bits_T_11 ? arr_38 : _GEN_3064; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3066 = 8'h27 == _io_out_bits_T_11 ? arr_39 : _GEN_3065; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3067 = 8'h28 == _io_out_bits_T_11 ? arr_40 : _GEN_3066; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3068 = 8'h29 == _io_out_bits_T_11 ? arr_41 : _GEN_3067; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3069 = 8'h2a == _io_out_bits_T_11 ? arr_42 : _GEN_3068; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3070 = 8'h2b == _io_out_bits_T_11 ? arr_43 : _GEN_3069; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3071 = 8'h2c == _io_out_bits_T_11 ? arr_44 : _GEN_3070; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3072 = 8'h2d == _io_out_bits_T_11 ? arr_45 : _GEN_3071; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3073 = 8'h2e == _io_out_bits_T_11 ? arr_46 : _GEN_3072; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3074 = 8'h2f == _io_out_bits_T_11 ? arr_47 : _GEN_3073; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3075 = 8'h30 == _io_out_bits_T_11 ? arr_48 : _GEN_3074; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3076 = 8'h31 == _io_out_bits_T_11 ? arr_49 : _GEN_3075; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3077 = 8'h32 == _io_out_bits_T_11 ? arr_50 : _GEN_3076; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3078 = 8'h33 == _io_out_bits_T_11 ? arr_51 : _GEN_3077; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3079 = 8'h34 == _io_out_bits_T_11 ? arr_52 : _GEN_3078; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3080 = 8'h35 == _io_out_bits_T_11 ? arr_53 : _GEN_3079; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3081 = 8'h36 == _io_out_bits_T_11 ? arr_54 : _GEN_3080; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3082 = 8'h37 == _io_out_bits_T_11 ? arr_55 : _GEN_3081; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3083 = 8'h38 == _io_out_bits_T_11 ? arr_56 : _GEN_3082; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3084 = 8'h39 == _io_out_bits_T_11 ? arr_57 : _GEN_3083; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3085 = 8'h3a == _io_out_bits_T_11 ? arr_58 : _GEN_3084; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3086 = 8'h3b == _io_out_bits_T_11 ? arr_59 : _GEN_3085; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3087 = 8'h3c == _io_out_bits_T_11 ? arr_60 : _GEN_3086; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3088 = 8'h3d == _io_out_bits_T_11 ? arr_61 : _GEN_3087; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3089 = 8'h3e == _io_out_bits_T_11 ? arr_62 : _GEN_3088; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3090 = 8'h3f == _io_out_bits_T_11 ? arr_63 : _GEN_3089; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3091 = 8'h40 == _io_out_bits_T_11 ? arr_64 : _GEN_3090; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3092 = 8'h41 == _io_out_bits_T_11 ? arr_65 : _GEN_3091; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3093 = 8'h42 == _io_out_bits_T_11 ? arr_66 : _GEN_3092; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3094 = 8'h43 == _io_out_bits_T_11 ? arr_67 : _GEN_3093; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3095 = 8'h44 == _io_out_bits_T_11 ? arr_68 : _GEN_3094; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3096 = 8'h45 == _io_out_bits_T_11 ? arr_69 : _GEN_3095; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3097 = 8'h46 == _io_out_bits_T_11 ? arr_70 : _GEN_3096; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3098 = 8'h47 == _io_out_bits_T_11 ? arr_71 : _GEN_3097; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3099 = 8'h48 == _io_out_bits_T_11 ? arr_72 : _GEN_3098; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3100 = 8'h49 == _io_out_bits_T_11 ? arr_73 : _GEN_3099; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3101 = 8'h4a == _io_out_bits_T_11 ? arr_74 : _GEN_3100; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3102 = 8'h4b == _io_out_bits_T_11 ? arr_75 : _GEN_3101; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3103 = 8'h4c == _io_out_bits_T_11 ? arr_76 : _GEN_3102; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3104 = 8'h4d == _io_out_bits_T_11 ? arr_77 : _GEN_3103; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3105 = 8'h4e == _io_out_bits_T_11 ? arr_78 : _GEN_3104; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3106 = 8'h4f == _io_out_bits_T_11 ? arr_79 : _GEN_3105; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3107 = 8'h50 == _io_out_bits_T_11 ? arr_80 : _GEN_3106; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3108 = 8'h51 == _io_out_bits_T_11 ? arr_81 : _GEN_3107; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3109 = 8'h52 == _io_out_bits_T_11 ? arr_82 : _GEN_3108; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3110 = 8'h53 == _io_out_bits_T_11 ? arr_83 : _GEN_3109; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3111 = 8'h54 == _io_out_bits_T_11 ? arr_84 : _GEN_3110; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3112 = 8'h55 == _io_out_bits_T_11 ? arr_85 : _GEN_3111; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3113 = 8'h56 == _io_out_bits_T_11 ? arr_86 : _GEN_3112; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3114 = 8'h57 == _io_out_bits_T_11 ? arr_87 : _GEN_3113; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3115 = 8'h58 == _io_out_bits_T_11 ? arr_88 : _GEN_3114; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3116 = 8'h59 == _io_out_bits_T_11 ? arr_89 : _GEN_3115; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3117 = 8'h5a == _io_out_bits_T_11 ? arr_90 : _GEN_3116; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3118 = 8'h5b == _io_out_bits_T_11 ? arr_91 : _GEN_3117; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3119 = 8'h5c == _io_out_bits_T_11 ? arr_92 : _GEN_3118; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3120 = 8'h5d == _io_out_bits_T_11 ? arr_93 : _GEN_3119; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3121 = 8'h5e == _io_out_bits_T_11 ? arr_94 : _GEN_3120; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3122 = 8'h5f == _io_out_bits_T_11 ? arr_95 : _GEN_3121; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3123 = 8'h60 == _io_out_bits_T_11 ? arr_96 : _GEN_3122; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3124 = 8'h61 == _io_out_bits_T_11 ? arr_97 : _GEN_3123; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3125 = 8'h62 == _io_out_bits_T_11 ? arr_98 : _GEN_3124; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3126 = 8'h63 == _io_out_bits_T_11 ? arr_99 : _GEN_3125; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3127 = 8'h64 == _io_out_bits_T_11 ? arr_100 : _GEN_3126; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3128 = 8'h65 == _io_out_bits_T_11 ? arr_101 : _GEN_3127; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3129 = 8'h66 == _io_out_bits_T_11 ? arr_102 : _GEN_3128; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3130 = 8'h67 == _io_out_bits_T_11 ? arr_103 : _GEN_3129; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3131 = 8'h68 == _io_out_bits_T_11 ? arr_104 : _GEN_3130; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3132 = 8'h69 == _io_out_bits_T_11 ? arr_105 : _GEN_3131; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3133 = 8'h6a == _io_out_bits_T_11 ? arr_106 : _GEN_3132; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3134 = 8'h6b == _io_out_bits_T_11 ? arr_107 : _GEN_3133; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3135 = 8'h6c == _io_out_bits_T_11 ? arr_108 : _GEN_3134; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3136 = 8'h6d == _io_out_bits_T_11 ? arr_109 : _GEN_3135; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3137 = 8'h6e == _io_out_bits_T_11 ? arr_110 : _GEN_3136; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3138 = 8'h6f == _io_out_bits_T_11 ? arr_111 : _GEN_3137; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3139 = 8'h70 == _io_out_bits_T_11 ? arr_112 : _GEN_3138; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3140 = 8'h71 == _io_out_bits_T_11 ? arr_113 : _GEN_3139; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3141 = 8'h72 == _io_out_bits_T_11 ? arr_114 : _GEN_3140; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3142 = 8'h73 == _io_out_bits_T_11 ? arr_115 : _GEN_3141; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3143 = 8'h74 == _io_out_bits_T_11 ? arr_116 : _GEN_3142; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3144 = 8'h75 == _io_out_bits_T_11 ? arr_117 : _GEN_3143; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3145 = 8'h76 == _io_out_bits_T_11 ? arr_118 : _GEN_3144; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3146 = 8'h77 == _io_out_bits_T_11 ? arr_119 : _GEN_3145; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3147 = 8'h78 == _io_out_bits_T_11 ? arr_120 : _GEN_3146; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3148 = 8'h79 == _io_out_bits_T_11 ? arr_121 : _GEN_3147; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3149 = 8'h7a == _io_out_bits_T_11 ? arr_122 : _GEN_3148; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3150 = 8'h7b == _io_out_bits_T_11 ? arr_123 : _GEN_3149; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3151 = 8'h7c == _io_out_bits_T_11 ? arr_124 : _GEN_3150; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3152 = 8'h7d == _io_out_bits_T_11 ? arr_125 : _GEN_3151; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3153 = 8'h7e == _io_out_bits_T_11 ? arr_126 : _GEN_3152; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3154 = 8'h7f == _io_out_bits_T_11 ? arr_127 : _GEN_3153; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3155 = 8'h80 == _io_out_bits_T_11 ? arr_128 : _GEN_3154; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3156 = 8'h81 == _io_out_bits_T_11 ? arr_129 : _GEN_3155; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3157 = 8'h82 == _io_out_bits_T_11 ? arr_130 : _GEN_3156; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3158 = 8'h83 == _io_out_bits_T_11 ? arr_131 : _GEN_3157; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3159 = 8'h84 == _io_out_bits_T_11 ? arr_132 : _GEN_3158; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3160 = 8'h85 == _io_out_bits_T_11 ? arr_133 : _GEN_3159; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3161 = 8'h86 == _io_out_bits_T_11 ? arr_134 : _GEN_3160; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3162 = 8'h87 == _io_out_bits_T_11 ? arr_135 : _GEN_3161; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3163 = 8'h88 == _io_out_bits_T_11 ? arr_136 : _GEN_3162; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3164 = 8'h89 == _io_out_bits_T_11 ? arr_137 : _GEN_3163; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3165 = 8'h8a == _io_out_bits_T_11 ? arr_138 : _GEN_3164; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3166 = 8'h8b == _io_out_bits_T_11 ? arr_139 : _GEN_3165; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3167 = 8'h8c == _io_out_bits_T_11 ? arr_140 : _GEN_3166; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3168 = 8'h8d == _io_out_bits_T_11 ? arr_141 : _GEN_3167; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3169 = 8'h8e == _io_out_bits_T_11 ? arr_142 : _GEN_3168; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3170 = 8'h8f == _io_out_bits_T_11 ? arr_143 : _GEN_3169; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3172 = 8'h1 == _io_out_bits_T_9 ? arr_1 : arr_0; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3173 = 8'h2 == _io_out_bits_T_9 ? arr_2 : _GEN_3172; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3174 = 8'h3 == _io_out_bits_T_9 ? arr_3 : _GEN_3173; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3175 = 8'h4 == _io_out_bits_T_9 ? arr_4 : _GEN_3174; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3176 = 8'h5 == _io_out_bits_T_9 ? arr_5 : _GEN_3175; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3177 = 8'h6 == _io_out_bits_T_9 ? arr_6 : _GEN_3176; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3178 = 8'h7 == _io_out_bits_T_9 ? arr_7 : _GEN_3177; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3179 = 8'h8 == _io_out_bits_T_9 ? arr_8 : _GEN_3178; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3180 = 8'h9 == _io_out_bits_T_9 ? arr_9 : _GEN_3179; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3181 = 8'ha == _io_out_bits_T_9 ? arr_10 : _GEN_3180; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3182 = 8'hb == _io_out_bits_T_9 ? arr_11 : _GEN_3181; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3183 = 8'hc == _io_out_bits_T_9 ? arr_12 : _GEN_3182; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3184 = 8'hd == _io_out_bits_T_9 ? arr_13 : _GEN_3183; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3185 = 8'he == _io_out_bits_T_9 ? arr_14 : _GEN_3184; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3186 = 8'hf == _io_out_bits_T_9 ? arr_15 : _GEN_3185; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3187 = 8'h10 == _io_out_bits_T_9 ? arr_16 : _GEN_3186; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3188 = 8'h11 == _io_out_bits_T_9 ? arr_17 : _GEN_3187; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3189 = 8'h12 == _io_out_bits_T_9 ? arr_18 : _GEN_3188; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3190 = 8'h13 == _io_out_bits_T_9 ? arr_19 : _GEN_3189; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3191 = 8'h14 == _io_out_bits_T_9 ? arr_20 : _GEN_3190; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3192 = 8'h15 == _io_out_bits_T_9 ? arr_21 : _GEN_3191; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3193 = 8'h16 == _io_out_bits_T_9 ? arr_22 : _GEN_3192; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3194 = 8'h17 == _io_out_bits_T_9 ? arr_23 : _GEN_3193; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3195 = 8'h18 == _io_out_bits_T_9 ? arr_24 : _GEN_3194; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3196 = 8'h19 == _io_out_bits_T_9 ? arr_25 : _GEN_3195; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3197 = 8'h1a == _io_out_bits_T_9 ? arr_26 : _GEN_3196; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3198 = 8'h1b == _io_out_bits_T_9 ? arr_27 : _GEN_3197; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3199 = 8'h1c == _io_out_bits_T_9 ? arr_28 : _GEN_3198; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3200 = 8'h1d == _io_out_bits_T_9 ? arr_29 : _GEN_3199; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3201 = 8'h1e == _io_out_bits_T_9 ? arr_30 : _GEN_3200; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3202 = 8'h1f == _io_out_bits_T_9 ? arr_31 : _GEN_3201; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3203 = 8'h20 == _io_out_bits_T_9 ? arr_32 : _GEN_3202; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3204 = 8'h21 == _io_out_bits_T_9 ? arr_33 : _GEN_3203; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3205 = 8'h22 == _io_out_bits_T_9 ? arr_34 : _GEN_3204; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3206 = 8'h23 == _io_out_bits_T_9 ? arr_35 : _GEN_3205; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3207 = 8'h24 == _io_out_bits_T_9 ? arr_36 : _GEN_3206; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3208 = 8'h25 == _io_out_bits_T_9 ? arr_37 : _GEN_3207; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3209 = 8'h26 == _io_out_bits_T_9 ? arr_38 : _GEN_3208; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3210 = 8'h27 == _io_out_bits_T_9 ? arr_39 : _GEN_3209; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3211 = 8'h28 == _io_out_bits_T_9 ? arr_40 : _GEN_3210; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3212 = 8'h29 == _io_out_bits_T_9 ? arr_41 : _GEN_3211; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3213 = 8'h2a == _io_out_bits_T_9 ? arr_42 : _GEN_3212; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3214 = 8'h2b == _io_out_bits_T_9 ? arr_43 : _GEN_3213; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3215 = 8'h2c == _io_out_bits_T_9 ? arr_44 : _GEN_3214; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3216 = 8'h2d == _io_out_bits_T_9 ? arr_45 : _GEN_3215; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3217 = 8'h2e == _io_out_bits_T_9 ? arr_46 : _GEN_3216; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3218 = 8'h2f == _io_out_bits_T_9 ? arr_47 : _GEN_3217; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3219 = 8'h30 == _io_out_bits_T_9 ? arr_48 : _GEN_3218; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3220 = 8'h31 == _io_out_bits_T_9 ? arr_49 : _GEN_3219; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3221 = 8'h32 == _io_out_bits_T_9 ? arr_50 : _GEN_3220; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3222 = 8'h33 == _io_out_bits_T_9 ? arr_51 : _GEN_3221; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3223 = 8'h34 == _io_out_bits_T_9 ? arr_52 : _GEN_3222; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3224 = 8'h35 == _io_out_bits_T_9 ? arr_53 : _GEN_3223; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3225 = 8'h36 == _io_out_bits_T_9 ? arr_54 : _GEN_3224; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3226 = 8'h37 == _io_out_bits_T_9 ? arr_55 : _GEN_3225; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3227 = 8'h38 == _io_out_bits_T_9 ? arr_56 : _GEN_3226; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3228 = 8'h39 == _io_out_bits_T_9 ? arr_57 : _GEN_3227; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3229 = 8'h3a == _io_out_bits_T_9 ? arr_58 : _GEN_3228; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3230 = 8'h3b == _io_out_bits_T_9 ? arr_59 : _GEN_3229; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3231 = 8'h3c == _io_out_bits_T_9 ? arr_60 : _GEN_3230; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3232 = 8'h3d == _io_out_bits_T_9 ? arr_61 : _GEN_3231; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3233 = 8'h3e == _io_out_bits_T_9 ? arr_62 : _GEN_3232; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3234 = 8'h3f == _io_out_bits_T_9 ? arr_63 : _GEN_3233; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3235 = 8'h40 == _io_out_bits_T_9 ? arr_64 : _GEN_3234; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3236 = 8'h41 == _io_out_bits_T_9 ? arr_65 : _GEN_3235; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3237 = 8'h42 == _io_out_bits_T_9 ? arr_66 : _GEN_3236; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3238 = 8'h43 == _io_out_bits_T_9 ? arr_67 : _GEN_3237; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3239 = 8'h44 == _io_out_bits_T_9 ? arr_68 : _GEN_3238; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3240 = 8'h45 == _io_out_bits_T_9 ? arr_69 : _GEN_3239; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3241 = 8'h46 == _io_out_bits_T_9 ? arr_70 : _GEN_3240; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3242 = 8'h47 == _io_out_bits_T_9 ? arr_71 : _GEN_3241; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3243 = 8'h48 == _io_out_bits_T_9 ? arr_72 : _GEN_3242; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3244 = 8'h49 == _io_out_bits_T_9 ? arr_73 : _GEN_3243; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3245 = 8'h4a == _io_out_bits_T_9 ? arr_74 : _GEN_3244; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3246 = 8'h4b == _io_out_bits_T_9 ? arr_75 : _GEN_3245; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3247 = 8'h4c == _io_out_bits_T_9 ? arr_76 : _GEN_3246; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3248 = 8'h4d == _io_out_bits_T_9 ? arr_77 : _GEN_3247; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3249 = 8'h4e == _io_out_bits_T_9 ? arr_78 : _GEN_3248; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3250 = 8'h4f == _io_out_bits_T_9 ? arr_79 : _GEN_3249; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3251 = 8'h50 == _io_out_bits_T_9 ? arr_80 : _GEN_3250; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3252 = 8'h51 == _io_out_bits_T_9 ? arr_81 : _GEN_3251; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3253 = 8'h52 == _io_out_bits_T_9 ? arr_82 : _GEN_3252; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3254 = 8'h53 == _io_out_bits_T_9 ? arr_83 : _GEN_3253; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3255 = 8'h54 == _io_out_bits_T_9 ? arr_84 : _GEN_3254; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3256 = 8'h55 == _io_out_bits_T_9 ? arr_85 : _GEN_3255; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3257 = 8'h56 == _io_out_bits_T_9 ? arr_86 : _GEN_3256; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3258 = 8'h57 == _io_out_bits_T_9 ? arr_87 : _GEN_3257; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3259 = 8'h58 == _io_out_bits_T_9 ? arr_88 : _GEN_3258; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3260 = 8'h59 == _io_out_bits_T_9 ? arr_89 : _GEN_3259; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3261 = 8'h5a == _io_out_bits_T_9 ? arr_90 : _GEN_3260; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3262 = 8'h5b == _io_out_bits_T_9 ? arr_91 : _GEN_3261; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3263 = 8'h5c == _io_out_bits_T_9 ? arr_92 : _GEN_3262; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3264 = 8'h5d == _io_out_bits_T_9 ? arr_93 : _GEN_3263; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3265 = 8'h5e == _io_out_bits_T_9 ? arr_94 : _GEN_3264; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3266 = 8'h5f == _io_out_bits_T_9 ? arr_95 : _GEN_3265; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3267 = 8'h60 == _io_out_bits_T_9 ? arr_96 : _GEN_3266; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3268 = 8'h61 == _io_out_bits_T_9 ? arr_97 : _GEN_3267; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3269 = 8'h62 == _io_out_bits_T_9 ? arr_98 : _GEN_3268; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3270 = 8'h63 == _io_out_bits_T_9 ? arr_99 : _GEN_3269; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3271 = 8'h64 == _io_out_bits_T_9 ? arr_100 : _GEN_3270; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3272 = 8'h65 == _io_out_bits_T_9 ? arr_101 : _GEN_3271; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3273 = 8'h66 == _io_out_bits_T_9 ? arr_102 : _GEN_3272; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3274 = 8'h67 == _io_out_bits_T_9 ? arr_103 : _GEN_3273; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3275 = 8'h68 == _io_out_bits_T_9 ? arr_104 : _GEN_3274; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3276 = 8'h69 == _io_out_bits_T_9 ? arr_105 : _GEN_3275; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3277 = 8'h6a == _io_out_bits_T_9 ? arr_106 : _GEN_3276; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3278 = 8'h6b == _io_out_bits_T_9 ? arr_107 : _GEN_3277; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3279 = 8'h6c == _io_out_bits_T_9 ? arr_108 : _GEN_3278; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3280 = 8'h6d == _io_out_bits_T_9 ? arr_109 : _GEN_3279; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3281 = 8'h6e == _io_out_bits_T_9 ? arr_110 : _GEN_3280; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3282 = 8'h6f == _io_out_bits_T_9 ? arr_111 : _GEN_3281; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3283 = 8'h70 == _io_out_bits_T_9 ? arr_112 : _GEN_3282; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3284 = 8'h71 == _io_out_bits_T_9 ? arr_113 : _GEN_3283; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3285 = 8'h72 == _io_out_bits_T_9 ? arr_114 : _GEN_3284; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3286 = 8'h73 == _io_out_bits_T_9 ? arr_115 : _GEN_3285; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3287 = 8'h74 == _io_out_bits_T_9 ? arr_116 : _GEN_3286; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3288 = 8'h75 == _io_out_bits_T_9 ? arr_117 : _GEN_3287; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3289 = 8'h76 == _io_out_bits_T_9 ? arr_118 : _GEN_3288; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3290 = 8'h77 == _io_out_bits_T_9 ? arr_119 : _GEN_3289; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3291 = 8'h78 == _io_out_bits_T_9 ? arr_120 : _GEN_3290; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3292 = 8'h79 == _io_out_bits_T_9 ? arr_121 : _GEN_3291; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3293 = 8'h7a == _io_out_bits_T_9 ? arr_122 : _GEN_3292; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3294 = 8'h7b == _io_out_bits_T_9 ? arr_123 : _GEN_3293; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3295 = 8'h7c == _io_out_bits_T_9 ? arr_124 : _GEN_3294; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3296 = 8'h7d == _io_out_bits_T_9 ? arr_125 : _GEN_3295; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3297 = 8'h7e == _io_out_bits_T_9 ? arr_126 : _GEN_3296; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3298 = 8'h7f == _io_out_bits_T_9 ? arr_127 : _GEN_3297; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3299 = 8'h80 == _io_out_bits_T_9 ? arr_128 : _GEN_3298; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3300 = 8'h81 == _io_out_bits_T_9 ? arr_129 : _GEN_3299; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3301 = 8'h82 == _io_out_bits_T_9 ? arr_130 : _GEN_3300; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3302 = 8'h83 == _io_out_bits_T_9 ? arr_131 : _GEN_3301; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3303 = 8'h84 == _io_out_bits_T_9 ? arr_132 : _GEN_3302; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3304 = 8'h85 == _io_out_bits_T_9 ? arr_133 : _GEN_3303; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3305 = 8'h86 == _io_out_bits_T_9 ? arr_134 : _GEN_3304; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3306 = 8'h87 == _io_out_bits_T_9 ? arr_135 : _GEN_3305; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3307 = 8'h88 == _io_out_bits_T_9 ? arr_136 : _GEN_3306; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3308 = 8'h89 == _io_out_bits_T_9 ? arr_137 : _GEN_3307; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3309 = 8'h8a == _io_out_bits_T_9 ? arr_138 : _GEN_3308; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3310 = 8'h8b == _io_out_bits_T_9 ? arr_139 : _GEN_3309; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3311 = 8'h8c == _io_out_bits_T_9 ? arr_140 : _GEN_3310; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3312 = 8'h8d == _io_out_bits_T_9 ? arr_141 : _GEN_3311; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3313 = 8'h8e == _io_out_bits_T_9 ? arr_142 : _GEN_3312; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3314 = 8'h8f == _io_out_bits_T_9 ? arr_143 : _GEN_3313; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3316 = 8'h1 == _io_out_bits_T_17 ? arr_1 : arr_0; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3317 = 8'h2 == _io_out_bits_T_17 ? arr_2 : _GEN_3316; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3318 = 8'h3 == _io_out_bits_T_17 ? arr_3 : _GEN_3317; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3319 = 8'h4 == _io_out_bits_T_17 ? arr_4 : _GEN_3318; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3320 = 8'h5 == _io_out_bits_T_17 ? arr_5 : _GEN_3319; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3321 = 8'h6 == _io_out_bits_T_17 ? arr_6 : _GEN_3320; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3322 = 8'h7 == _io_out_bits_T_17 ? arr_7 : _GEN_3321; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3323 = 8'h8 == _io_out_bits_T_17 ? arr_8 : _GEN_3322; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3324 = 8'h9 == _io_out_bits_T_17 ? arr_9 : _GEN_3323; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3325 = 8'ha == _io_out_bits_T_17 ? arr_10 : _GEN_3324; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3326 = 8'hb == _io_out_bits_T_17 ? arr_11 : _GEN_3325; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3327 = 8'hc == _io_out_bits_T_17 ? arr_12 : _GEN_3326; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3328 = 8'hd == _io_out_bits_T_17 ? arr_13 : _GEN_3327; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3329 = 8'he == _io_out_bits_T_17 ? arr_14 : _GEN_3328; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3330 = 8'hf == _io_out_bits_T_17 ? arr_15 : _GEN_3329; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3331 = 8'h10 == _io_out_bits_T_17 ? arr_16 : _GEN_3330; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3332 = 8'h11 == _io_out_bits_T_17 ? arr_17 : _GEN_3331; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3333 = 8'h12 == _io_out_bits_T_17 ? arr_18 : _GEN_3332; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3334 = 8'h13 == _io_out_bits_T_17 ? arr_19 : _GEN_3333; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3335 = 8'h14 == _io_out_bits_T_17 ? arr_20 : _GEN_3334; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3336 = 8'h15 == _io_out_bits_T_17 ? arr_21 : _GEN_3335; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3337 = 8'h16 == _io_out_bits_T_17 ? arr_22 : _GEN_3336; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3338 = 8'h17 == _io_out_bits_T_17 ? arr_23 : _GEN_3337; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3339 = 8'h18 == _io_out_bits_T_17 ? arr_24 : _GEN_3338; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3340 = 8'h19 == _io_out_bits_T_17 ? arr_25 : _GEN_3339; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3341 = 8'h1a == _io_out_bits_T_17 ? arr_26 : _GEN_3340; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3342 = 8'h1b == _io_out_bits_T_17 ? arr_27 : _GEN_3341; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3343 = 8'h1c == _io_out_bits_T_17 ? arr_28 : _GEN_3342; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3344 = 8'h1d == _io_out_bits_T_17 ? arr_29 : _GEN_3343; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3345 = 8'h1e == _io_out_bits_T_17 ? arr_30 : _GEN_3344; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3346 = 8'h1f == _io_out_bits_T_17 ? arr_31 : _GEN_3345; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3347 = 8'h20 == _io_out_bits_T_17 ? arr_32 : _GEN_3346; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3348 = 8'h21 == _io_out_bits_T_17 ? arr_33 : _GEN_3347; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3349 = 8'h22 == _io_out_bits_T_17 ? arr_34 : _GEN_3348; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3350 = 8'h23 == _io_out_bits_T_17 ? arr_35 : _GEN_3349; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3351 = 8'h24 == _io_out_bits_T_17 ? arr_36 : _GEN_3350; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3352 = 8'h25 == _io_out_bits_T_17 ? arr_37 : _GEN_3351; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3353 = 8'h26 == _io_out_bits_T_17 ? arr_38 : _GEN_3352; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3354 = 8'h27 == _io_out_bits_T_17 ? arr_39 : _GEN_3353; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3355 = 8'h28 == _io_out_bits_T_17 ? arr_40 : _GEN_3354; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3356 = 8'h29 == _io_out_bits_T_17 ? arr_41 : _GEN_3355; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3357 = 8'h2a == _io_out_bits_T_17 ? arr_42 : _GEN_3356; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3358 = 8'h2b == _io_out_bits_T_17 ? arr_43 : _GEN_3357; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3359 = 8'h2c == _io_out_bits_T_17 ? arr_44 : _GEN_3358; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3360 = 8'h2d == _io_out_bits_T_17 ? arr_45 : _GEN_3359; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3361 = 8'h2e == _io_out_bits_T_17 ? arr_46 : _GEN_3360; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3362 = 8'h2f == _io_out_bits_T_17 ? arr_47 : _GEN_3361; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3363 = 8'h30 == _io_out_bits_T_17 ? arr_48 : _GEN_3362; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3364 = 8'h31 == _io_out_bits_T_17 ? arr_49 : _GEN_3363; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3365 = 8'h32 == _io_out_bits_T_17 ? arr_50 : _GEN_3364; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3366 = 8'h33 == _io_out_bits_T_17 ? arr_51 : _GEN_3365; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3367 = 8'h34 == _io_out_bits_T_17 ? arr_52 : _GEN_3366; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3368 = 8'h35 == _io_out_bits_T_17 ? arr_53 : _GEN_3367; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3369 = 8'h36 == _io_out_bits_T_17 ? arr_54 : _GEN_3368; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3370 = 8'h37 == _io_out_bits_T_17 ? arr_55 : _GEN_3369; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3371 = 8'h38 == _io_out_bits_T_17 ? arr_56 : _GEN_3370; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3372 = 8'h39 == _io_out_bits_T_17 ? arr_57 : _GEN_3371; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3373 = 8'h3a == _io_out_bits_T_17 ? arr_58 : _GEN_3372; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3374 = 8'h3b == _io_out_bits_T_17 ? arr_59 : _GEN_3373; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3375 = 8'h3c == _io_out_bits_T_17 ? arr_60 : _GEN_3374; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3376 = 8'h3d == _io_out_bits_T_17 ? arr_61 : _GEN_3375; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3377 = 8'h3e == _io_out_bits_T_17 ? arr_62 : _GEN_3376; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3378 = 8'h3f == _io_out_bits_T_17 ? arr_63 : _GEN_3377; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3379 = 8'h40 == _io_out_bits_T_17 ? arr_64 : _GEN_3378; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3380 = 8'h41 == _io_out_bits_T_17 ? arr_65 : _GEN_3379; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3381 = 8'h42 == _io_out_bits_T_17 ? arr_66 : _GEN_3380; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3382 = 8'h43 == _io_out_bits_T_17 ? arr_67 : _GEN_3381; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3383 = 8'h44 == _io_out_bits_T_17 ? arr_68 : _GEN_3382; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3384 = 8'h45 == _io_out_bits_T_17 ? arr_69 : _GEN_3383; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3385 = 8'h46 == _io_out_bits_T_17 ? arr_70 : _GEN_3384; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3386 = 8'h47 == _io_out_bits_T_17 ? arr_71 : _GEN_3385; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3387 = 8'h48 == _io_out_bits_T_17 ? arr_72 : _GEN_3386; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3388 = 8'h49 == _io_out_bits_T_17 ? arr_73 : _GEN_3387; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3389 = 8'h4a == _io_out_bits_T_17 ? arr_74 : _GEN_3388; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3390 = 8'h4b == _io_out_bits_T_17 ? arr_75 : _GEN_3389; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3391 = 8'h4c == _io_out_bits_T_17 ? arr_76 : _GEN_3390; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3392 = 8'h4d == _io_out_bits_T_17 ? arr_77 : _GEN_3391; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3393 = 8'h4e == _io_out_bits_T_17 ? arr_78 : _GEN_3392; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3394 = 8'h4f == _io_out_bits_T_17 ? arr_79 : _GEN_3393; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3395 = 8'h50 == _io_out_bits_T_17 ? arr_80 : _GEN_3394; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3396 = 8'h51 == _io_out_bits_T_17 ? arr_81 : _GEN_3395; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3397 = 8'h52 == _io_out_bits_T_17 ? arr_82 : _GEN_3396; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3398 = 8'h53 == _io_out_bits_T_17 ? arr_83 : _GEN_3397; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3399 = 8'h54 == _io_out_bits_T_17 ? arr_84 : _GEN_3398; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3400 = 8'h55 == _io_out_bits_T_17 ? arr_85 : _GEN_3399; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3401 = 8'h56 == _io_out_bits_T_17 ? arr_86 : _GEN_3400; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3402 = 8'h57 == _io_out_bits_T_17 ? arr_87 : _GEN_3401; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3403 = 8'h58 == _io_out_bits_T_17 ? arr_88 : _GEN_3402; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3404 = 8'h59 == _io_out_bits_T_17 ? arr_89 : _GEN_3403; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3405 = 8'h5a == _io_out_bits_T_17 ? arr_90 : _GEN_3404; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3406 = 8'h5b == _io_out_bits_T_17 ? arr_91 : _GEN_3405; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3407 = 8'h5c == _io_out_bits_T_17 ? arr_92 : _GEN_3406; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3408 = 8'h5d == _io_out_bits_T_17 ? arr_93 : _GEN_3407; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3409 = 8'h5e == _io_out_bits_T_17 ? arr_94 : _GEN_3408; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3410 = 8'h5f == _io_out_bits_T_17 ? arr_95 : _GEN_3409; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3411 = 8'h60 == _io_out_bits_T_17 ? arr_96 : _GEN_3410; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3412 = 8'h61 == _io_out_bits_T_17 ? arr_97 : _GEN_3411; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3413 = 8'h62 == _io_out_bits_T_17 ? arr_98 : _GEN_3412; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3414 = 8'h63 == _io_out_bits_T_17 ? arr_99 : _GEN_3413; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3415 = 8'h64 == _io_out_bits_T_17 ? arr_100 : _GEN_3414; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3416 = 8'h65 == _io_out_bits_T_17 ? arr_101 : _GEN_3415; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3417 = 8'h66 == _io_out_bits_T_17 ? arr_102 : _GEN_3416; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3418 = 8'h67 == _io_out_bits_T_17 ? arr_103 : _GEN_3417; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3419 = 8'h68 == _io_out_bits_T_17 ? arr_104 : _GEN_3418; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3420 = 8'h69 == _io_out_bits_T_17 ? arr_105 : _GEN_3419; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3421 = 8'h6a == _io_out_bits_T_17 ? arr_106 : _GEN_3420; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3422 = 8'h6b == _io_out_bits_T_17 ? arr_107 : _GEN_3421; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3423 = 8'h6c == _io_out_bits_T_17 ? arr_108 : _GEN_3422; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3424 = 8'h6d == _io_out_bits_T_17 ? arr_109 : _GEN_3423; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3425 = 8'h6e == _io_out_bits_T_17 ? arr_110 : _GEN_3424; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3426 = 8'h6f == _io_out_bits_T_17 ? arr_111 : _GEN_3425; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3427 = 8'h70 == _io_out_bits_T_17 ? arr_112 : _GEN_3426; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3428 = 8'h71 == _io_out_bits_T_17 ? arr_113 : _GEN_3427; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3429 = 8'h72 == _io_out_bits_T_17 ? arr_114 : _GEN_3428; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3430 = 8'h73 == _io_out_bits_T_17 ? arr_115 : _GEN_3429; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3431 = 8'h74 == _io_out_bits_T_17 ? arr_116 : _GEN_3430; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3432 = 8'h75 == _io_out_bits_T_17 ? arr_117 : _GEN_3431; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3433 = 8'h76 == _io_out_bits_T_17 ? arr_118 : _GEN_3432; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3434 = 8'h77 == _io_out_bits_T_17 ? arr_119 : _GEN_3433; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3435 = 8'h78 == _io_out_bits_T_17 ? arr_120 : _GEN_3434; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3436 = 8'h79 == _io_out_bits_T_17 ? arr_121 : _GEN_3435; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3437 = 8'h7a == _io_out_bits_T_17 ? arr_122 : _GEN_3436; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3438 = 8'h7b == _io_out_bits_T_17 ? arr_123 : _GEN_3437; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3439 = 8'h7c == _io_out_bits_T_17 ? arr_124 : _GEN_3438; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3440 = 8'h7d == _io_out_bits_T_17 ? arr_125 : _GEN_3439; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3441 = 8'h7e == _io_out_bits_T_17 ? arr_126 : _GEN_3440; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3442 = 8'h7f == _io_out_bits_T_17 ? arr_127 : _GEN_3441; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3443 = 8'h80 == _io_out_bits_T_17 ? arr_128 : _GEN_3442; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3444 = 8'h81 == _io_out_bits_T_17 ? arr_129 : _GEN_3443; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3445 = 8'h82 == _io_out_bits_T_17 ? arr_130 : _GEN_3444; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3446 = 8'h83 == _io_out_bits_T_17 ? arr_131 : _GEN_3445; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3447 = 8'h84 == _io_out_bits_T_17 ? arr_132 : _GEN_3446; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3448 = 8'h85 == _io_out_bits_T_17 ? arr_133 : _GEN_3447; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3449 = 8'h86 == _io_out_bits_T_17 ? arr_134 : _GEN_3448; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3450 = 8'h87 == _io_out_bits_T_17 ? arr_135 : _GEN_3449; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3451 = 8'h88 == _io_out_bits_T_17 ? arr_136 : _GEN_3450; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3452 = 8'h89 == _io_out_bits_T_17 ? arr_137 : _GEN_3451; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3453 = 8'h8a == _io_out_bits_T_17 ? arr_138 : _GEN_3452; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3454 = 8'h8b == _io_out_bits_T_17 ? arr_139 : _GEN_3453; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3455 = 8'h8c == _io_out_bits_T_17 ? arr_140 : _GEN_3454; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3456 = 8'h8d == _io_out_bits_T_17 ? arr_141 : _GEN_3455; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3457 = 8'h8e == _io_out_bits_T_17 ? arr_142 : _GEN_3456; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3458 = 8'h8f == _io_out_bits_T_17 ? arr_143 : _GEN_3457; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3460 = 8'h1 == _io_out_bits_T_15 ? arr_1 : arr_0; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3461 = 8'h2 == _io_out_bits_T_15 ? arr_2 : _GEN_3460; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3462 = 8'h3 == _io_out_bits_T_15 ? arr_3 : _GEN_3461; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3463 = 8'h4 == _io_out_bits_T_15 ? arr_4 : _GEN_3462; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3464 = 8'h5 == _io_out_bits_T_15 ? arr_5 : _GEN_3463; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3465 = 8'h6 == _io_out_bits_T_15 ? arr_6 : _GEN_3464; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3466 = 8'h7 == _io_out_bits_T_15 ? arr_7 : _GEN_3465; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3467 = 8'h8 == _io_out_bits_T_15 ? arr_8 : _GEN_3466; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3468 = 8'h9 == _io_out_bits_T_15 ? arr_9 : _GEN_3467; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3469 = 8'ha == _io_out_bits_T_15 ? arr_10 : _GEN_3468; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3470 = 8'hb == _io_out_bits_T_15 ? arr_11 : _GEN_3469; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3471 = 8'hc == _io_out_bits_T_15 ? arr_12 : _GEN_3470; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3472 = 8'hd == _io_out_bits_T_15 ? arr_13 : _GEN_3471; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3473 = 8'he == _io_out_bits_T_15 ? arr_14 : _GEN_3472; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3474 = 8'hf == _io_out_bits_T_15 ? arr_15 : _GEN_3473; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3475 = 8'h10 == _io_out_bits_T_15 ? arr_16 : _GEN_3474; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3476 = 8'h11 == _io_out_bits_T_15 ? arr_17 : _GEN_3475; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3477 = 8'h12 == _io_out_bits_T_15 ? arr_18 : _GEN_3476; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3478 = 8'h13 == _io_out_bits_T_15 ? arr_19 : _GEN_3477; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3479 = 8'h14 == _io_out_bits_T_15 ? arr_20 : _GEN_3478; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3480 = 8'h15 == _io_out_bits_T_15 ? arr_21 : _GEN_3479; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3481 = 8'h16 == _io_out_bits_T_15 ? arr_22 : _GEN_3480; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3482 = 8'h17 == _io_out_bits_T_15 ? arr_23 : _GEN_3481; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3483 = 8'h18 == _io_out_bits_T_15 ? arr_24 : _GEN_3482; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3484 = 8'h19 == _io_out_bits_T_15 ? arr_25 : _GEN_3483; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3485 = 8'h1a == _io_out_bits_T_15 ? arr_26 : _GEN_3484; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3486 = 8'h1b == _io_out_bits_T_15 ? arr_27 : _GEN_3485; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3487 = 8'h1c == _io_out_bits_T_15 ? arr_28 : _GEN_3486; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3488 = 8'h1d == _io_out_bits_T_15 ? arr_29 : _GEN_3487; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3489 = 8'h1e == _io_out_bits_T_15 ? arr_30 : _GEN_3488; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3490 = 8'h1f == _io_out_bits_T_15 ? arr_31 : _GEN_3489; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3491 = 8'h20 == _io_out_bits_T_15 ? arr_32 : _GEN_3490; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3492 = 8'h21 == _io_out_bits_T_15 ? arr_33 : _GEN_3491; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3493 = 8'h22 == _io_out_bits_T_15 ? arr_34 : _GEN_3492; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3494 = 8'h23 == _io_out_bits_T_15 ? arr_35 : _GEN_3493; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3495 = 8'h24 == _io_out_bits_T_15 ? arr_36 : _GEN_3494; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3496 = 8'h25 == _io_out_bits_T_15 ? arr_37 : _GEN_3495; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3497 = 8'h26 == _io_out_bits_T_15 ? arr_38 : _GEN_3496; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3498 = 8'h27 == _io_out_bits_T_15 ? arr_39 : _GEN_3497; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3499 = 8'h28 == _io_out_bits_T_15 ? arr_40 : _GEN_3498; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3500 = 8'h29 == _io_out_bits_T_15 ? arr_41 : _GEN_3499; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3501 = 8'h2a == _io_out_bits_T_15 ? arr_42 : _GEN_3500; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3502 = 8'h2b == _io_out_bits_T_15 ? arr_43 : _GEN_3501; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3503 = 8'h2c == _io_out_bits_T_15 ? arr_44 : _GEN_3502; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3504 = 8'h2d == _io_out_bits_T_15 ? arr_45 : _GEN_3503; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3505 = 8'h2e == _io_out_bits_T_15 ? arr_46 : _GEN_3504; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3506 = 8'h2f == _io_out_bits_T_15 ? arr_47 : _GEN_3505; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3507 = 8'h30 == _io_out_bits_T_15 ? arr_48 : _GEN_3506; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3508 = 8'h31 == _io_out_bits_T_15 ? arr_49 : _GEN_3507; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3509 = 8'h32 == _io_out_bits_T_15 ? arr_50 : _GEN_3508; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3510 = 8'h33 == _io_out_bits_T_15 ? arr_51 : _GEN_3509; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3511 = 8'h34 == _io_out_bits_T_15 ? arr_52 : _GEN_3510; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3512 = 8'h35 == _io_out_bits_T_15 ? arr_53 : _GEN_3511; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3513 = 8'h36 == _io_out_bits_T_15 ? arr_54 : _GEN_3512; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3514 = 8'h37 == _io_out_bits_T_15 ? arr_55 : _GEN_3513; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3515 = 8'h38 == _io_out_bits_T_15 ? arr_56 : _GEN_3514; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3516 = 8'h39 == _io_out_bits_T_15 ? arr_57 : _GEN_3515; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3517 = 8'h3a == _io_out_bits_T_15 ? arr_58 : _GEN_3516; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3518 = 8'h3b == _io_out_bits_T_15 ? arr_59 : _GEN_3517; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3519 = 8'h3c == _io_out_bits_T_15 ? arr_60 : _GEN_3518; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3520 = 8'h3d == _io_out_bits_T_15 ? arr_61 : _GEN_3519; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3521 = 8'h3e == _io_out_bits_T_15 ? arr_62 : _GEN_3520; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3522 = 8'h3f == _io_out_bits_T_15 ? arr_63 : _GEN_3521; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3523 = 8'h40 == _io_out_bits_T_15 ? arr_64 : _GEN_3522; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3524 = 8'h41 == _io_out_bits_T_15 ? arr_65 : _GEN_3523; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3525 = 8'h42 == _io_out_bits_T_15 ? arr_66 : _GEN_3524; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3526 = 8'h43 == _io_out_bits_T_15 ? arr_67 : _GEN_3525; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3527 = 8'h44 == _io_out_bits_T_15 ? arr_68 : _GEN_3526; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3528 = 8'h45 == _io_out_bits_T_15 ? arr_69 : _GEN_3527; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3529 = 8'h46 == _io_out_bits_T_15 ? arr_70 : _GEN_3528; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3530 = 8'h47 == _io_out_bits_T_15 ? arr_71 : _GEN_3529; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3531 = 8'h48 == _io_out_bits_T_15 ? arr_72 : _GEN_3530; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3532 = 8'h49 == _io_out_bits_T_15 ? arr_73 : _GEN_3531; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3533 = 8'h4a == _io_out_bits_T_15 ? arr_74 : _GEN_3532; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3534 = 8'h4b == _io_out_bits_T_15 ? arr_75 : _GEN_3533; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3535 = 8'h4c == _io_out_bits_T_15 ? arr_76 : _GEN_3534; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3536 = 8'h4d == _io_out_bits_T_15 ? arr_77 : _GEN_3535; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3537 = 8'h4e == _io_out_bits_T_15 ? arr_78 : _GEN_3536; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3538 = 8'h4f == _io_out_bits_T_15 ? arr_79 : _GEN_3537; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3539 = 8'h50 == _io_out_bits_T_15 ? arr_80 : _GEN_3538; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3540 = 8'h51 == _io_out_bits_T_15 ? arr_81 : _GEN_3539; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3541 = 8'h52 == _io_out_bits_T_15 ? arr_82 : _GEN_3540; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3542 = 8'h53 == _io_out_bits_T_15 ? arr_83 : _GEN_3541; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3543 = 8'h54 == _io_out_bits_T_15 ? arr_84 : _GEN_3542; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3544 = 8'h55 == _io_out_bits_T_15 ? arr_85 : _GEN_3543; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3545 = 8'h56 == _io_out_bits_T_15 ? arr_86 : _GEN_3544; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3546 = 8'h57 == _io_out_bits_T_15 ? arr_87 : _GEN_3545; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3547 = 8'h58 == _io_out_bits_T_15 ? arr_88 : _GEN_3546; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3548 = 8'h59 == _io_out_bits_T_15 ? arr_89 : _GEN_3547; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3549 = 8'h5a == _io_out_bits_T_15 ? arr_90 : _GEN_3548; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3550 = 8'h5b == _io_out_bits_T_15 ? arr_91 : _GEN_3549; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3551 = 8'h5c == _io_out_bits_T_15 ? arr_92 : _GEN_3550; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3552 = 8'h5d == _io_out_bits_T_15 ? arr_93 : _GEN_3551; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3553 = 8'h5e == _io_out_bits_T_15 ? arr_94 : _GEN_3552; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3554 = 8'h5f == _io_out_bits_T_15 ? arr_95 : _GEN_3553; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3555 = 8'h60 == _io_out_bits_T_15 ? arr_96 : _GEN_3554; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3556 = 8'h61 == _io_out_bits_T_15 ? arr_97 : _GEN_3555; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3557 = 8'h62 == _io_out_bits_T_15 ? arr_98 : _GEN_3556; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3558 = 8'h63 == _io_out_bits_T_15 ? arr_99 : _GEN_3557; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3559 = 8'h64 == _io_out_bits_T_15 ? arr_100 : _GEN_3558; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3560 = 8'h65 == _io_out_bits_T_15 ? arr_101 : _GEN_3559; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3561 = 8'h66 == _io_out_bits_T_15 ? arr_102 : _GEN_3560; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3562 = 8'h67 == _io_out_bits_T_15 ? arr_103 : _GEN_3561; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3563 = 8'h68 == _io_out_bits_T_15 ? arr_104 : _GEN_3562; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3564 = 8'h69 == _io_out_bits_T_15 ? arr_105 : _GEN_3563; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3565 = 8'h6a == _io_out_bits_T_15 ? arr_106 : _GEN_3564; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3566 = 8'h6b == _io_out_bits_T_15 ? arr_107 : _GEN_3565; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3567 = 8'h6c == _io_out_bits_T_15 ? arr_108 : _GEN_3566; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3568 = 8'h6d == _io_out_bits_T_15 ? arr_109 : _GEN_3567; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3569 = 8'h6e == _io_out_bits_T_15 ? arr_110 : _GEN_3568; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3570 = 8'h6f == _io_out_bits_T_15 ? arr_111 : _GEN_3569; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3571 = 8'h70 == _io_out_bits_T_15 ? arr_112 : _GEN_3570; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3572 = 8'h71 == _io_out_bits_T_15 ? arr_113 : _GEN_3571; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3573 = 8'h72 == _io_out_bits_T_15 ? arr_114 : _GEN_3572; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3574 = 8'h73 == _io_out_bits_T_15 ? arr_115 : _GEN_3573; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3575 = 8'h74 == _io_out_bits_T_15 ? arr_116 : _GEN_3574; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3576 = 8'h75 == _io_out_bits_T_15 ? arr_117 : _GEN_3575; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3577 = 8'h76 == _io_out_bits_T_15 ? arr_118 : _GEN_3576; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3578 = 8'h77 == _io_out_bits_T_15 ? arr_119 : _GEN_3577; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3579 = 8'h78 == _io_out_bits_T_15 ? arr_120 : _GEN_3578; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3580 = 8'h79 == _io_out_bits_T_15 ? arr_121 : _GEN_3579; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3581 = 8'h7a == _io_out_bits_T_15 ? arr_122 : _GEN_3580; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3582 = 8'h7b == _io_out_bits_T_15 ? arr_123 : _GEN_3581; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3583 = 8'h7c == _io_out_bits_T_15 ? arr_124 : _GEN_3582; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3584 = 8'h7d == _io_out_bits_T_15 ? arr_125 : _GEN_3583; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3585 = 8'h7e == _io_out_bits_T_15 ? arr_126 : _GEN_3584; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3586 = 8'h7f == _io_out_bits_T_15 ? arr_127 : _GEN_3585; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3587 = 8'h80 == _io_out_bits_T_15 ? arr_128 : _GEN_3586; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3588 = 8'h81 == _io_out_bits_T_15 ? arr_129 : _GEN_3587; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3589 = 8'h82 == _io_out_bits_T_15 ? arr_130 : _GEN_3588; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3590 = 8'h83 == _io_out_bits_T_15 ? arr_131 : _GEN_3589; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3591 = 8'h84 == _io_out_bits_T_15 ? arr_132 : _GEN_3590; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3592 = 8'h85 == _io_out_bits_T_15 ? arr_133 : _GEN_3591; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3593 = 8'h86 == _io_out_bits_T_15 ? arr_134 : _GEN_3592; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3594 = 8'h87 == _io_out_bits_T_15 ? arr_135 : _GEN_3593; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3595 = 8'h88 == _io_out_bits_T_15 ? arr_136 : _GEN_3594; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3596 = 8'h89 == _io_out_bits_T_15 ? arr_137 : _GEN_3595; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3597 = 8'h8a == _io_out_bits_T_15 ? arr_138 : _GEN_3596; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3598 = 8'h8b == _io_out_bits_T_15 ? arr_139 : _GEN_3597; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3599 = 8'h8c == _io_out_bits_T_15 ? arr_140 : _GEN_3598; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3600 = 8'h8d == _io_out_bits_T_15 ? arr_141 : _GEN_3599; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3601 = 8'h8e == _io_out_bits_T_15 ? arr_142 : _GEN_3600; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3602 = 8'h8f == _io_out_bits_T_15 ? arr_143 : _GEN_3601; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3604 = 8'h1 == _io_out_bits_T_13 ? arr_1 : arr_0; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3605 = 8'h2 == _io_out_bits_T_13 ? arr_2 : _GEN_3604; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3606 = 8'h3 == _io_out_bits_T_13 ? arr_3 : _GEN_3605; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3607 = 8'h4 == _io_out_bits_T_13 ? arr_4 : _GEN_3606; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3608 = 8'h5 == _io_out_bits_T_13 ? arr_5 : _GEN_3607; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3609 = 8'h6 == _io_out_bits_T_13 ? arr_6 : _GEN_3608; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3610 = 8'h7 == _io_out_bits_T_13 ? arr_7 : _GEN_3609; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3611 = 8'h8 == _io_out_bits_T_13 ? arr_8 : _GEN_3610; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3612 = 8'h9 == _io_out_bits_T_13 ? arr_9 : _GEN_3611; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3613 = 8'ha == _io_out_bits_T_13 ? arr_10 : _GEN_3612; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3614 = 8'hb == _io_out_bits_T_13 ? arr_11 : _GEN_3613; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3615 = 8'hc == _io_out_bits_T_13 ? arr_12 : _GEN_3614; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3616 = 8'hd == _io_out_bits_T_13 ? arr_13 : _GEN_3615; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3617 = 8'he == _io_out_bits_T_13 ? arr_14 : _GEN_3616; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3618 = 8'hf == _io_out_bits_T_13 ? arr_15 : _GEN_3617; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3619 = 8'h10 == _io_out_bits_T_13 ? arr_16 : _GEN_3618; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3620 = 8'h11 == _io_out_bits_T_13 ? arr_17 : _GEN_3619; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3621 = 8'h12 == _io_out_bits_T_13 ? arr_18 : _GEN_3620; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3622 = 8'h13 == _io_out_bits_T_13 ? arr_19 : _GEN_3621; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3623 = 8'h14 == _io_out_bits_T_13 ? arr_20 : _GEN_3622; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3624 = 8'h15 == _io_out_bits_T_13 ? arr_21 : _GEN_3623; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3625 = 8'h16 == _io_out_bits_T_13 ? arr_22 : _GEN_3624; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3626 = 8'h17 == _io_out_bits_T_13 ? arr_23 : _GEN_3625; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3627 = 8'h18 == _io_out_bits_T_13 ? arr_24 : _GEN_3626; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3628 = 8'h19 == _io_out_bits_T_13 ? arr_25 : _GEN_3627; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3629 = 8'h1a == _io_out_bits_T_13 ? arr_26 : _GEN_3628; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3630 = 8'h1b == _io_out_bits_T_13 ? arr_27 : _GEN_3629; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3631 = 8'h1c == _io_out_bits_T_13 ? arr_28 : _GEN_3630; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3632 = 8'h1d == _io_out_bits_T_13 ? arr_29 : _GEN_3631; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3633 = 8'h1e == _io_out_bits_T_13 ? arr_30 : _GEN_3632; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3634 = 8'h1f == _io_out_bits_T_13 ? arr_31 : _GEN_3633; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3635 = 8'h20 == _io_out_bits_T_13 ? arr_32 : _GEN_3634; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3636 = 8'h21 == _io_out_bits_T_13 ? arr_33 : _GEN_3635; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3637 = 8'h22 == _io_out_bits_T_13 ? arr_34 : _GEN_3636; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3638 = 8'h23 == _io_out_bits_T_13 ? arr_35 : _GEN_3637; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3639 = 8'h24 == _io_out_bits_T_13 ? arr_36 : _GEN_3638; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3640 = 8'h25 == _io_out_bits_T_13 ? arr_37 : _GEN_3639; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3641 = 8'h26 == _io_out_bits_T_13 ? arr_38 : _GEN_3640; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3642 = 8'h27 == _io_out_bits_T_13 ? arr_39 : _GEN_3641; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3643 = 8'h28 == _io_out_bits_T_13 ? arr_40 : _GEN_3642; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3644 = 8'h29 == _io_out_bits_T_13 ? arr_41 : _GEN_3643; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3645 = 8'h2a == _io_out_bits_T_13 ? arr_42 : _GEN_3644; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3646 = 8'h2b == _io_out_bits_T_13 ? arr_43 : _GEN_3645; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3647 = 8'h2c == _io_out_bits_T_13 ? arr_44 : _GEN_3646; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3648 = 8'h2d == _io_out_bits_T_13 ? arr_45 : _GEN_3647; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3649 = 8'h2e == _io_out_bits_T_13 ? arr_46 : _GEN_3648; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3650 = 8'h2f == _io_out_bits_T_13 ? arr_47 : _GEN_3649; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3651 = 8'h30 == _io_out_bits_T_13 ? arr_48 : _GEN_3650; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3652 = 8'h31 == _io_out_bits_T_13 ? arr_49 : _GEN_3651; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3653 = 8'h32 == _io_out_bits_T_13 ? arr_50 : _GEN_3652; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3654 = 8'h33 == _io_out_bits_T_13 ? arr_51 : _GEN_3653; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3655 = 8'h34 == _io_out_bits_T_13 ? arr_52 : _GEN_3654; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3656 = 8'h35 == _io_out_bits_T_13 ? arr_53 : _GEN_3655; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3657 = 8'h36 == _io_out_bits_T_13 ? arr_54 : _GEN_3656; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3658 = 8'h37 == _io_out_bits_T_13 ? arr_55 : _GEN_3657; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3659 = 8'h38 == _io_out_bits_T_13 ? arr_56 : _GEN_3658; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3660 = 8'h39 == _io_out_bits_T_13 ? arr_57 : _GEN_3659; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3661 = 8'h3a == _io_out_bits_T_13 ? arr_58 : _GEN_3660; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3662 = 8'h3b == _io_out_bits_T_13 ? arr_59 : _GEN_3661; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3663 = 8'h3c == _io_out_bits_T_13 ? arr_60 : _GEN_3662; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3664 = 8'h3d == _io_out_bits_T_13 ? arr_61 : _GEN_3663; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3665 = 8'h3e == _io_out_bits_T_13 ? arr_62 : _GEN_3664; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3666 = 8'h3f == _io_out_bits_T_13 ? arr_63 : _GEN_3665; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3667 = 8'h40 == _io_out_bits_T_13 ? arr_64 : _GEN_3666; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3668 = 8'h41 == _io_out_bits_T_13 ? arr_65 : _GEN_3667; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3669 = 8'h42 == _io_out_bits_T_13 ? arr_66 : _GEN_3668; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3670 = 8'h43 == _io_out_bits_T_13 ? arr_67 : _GEN_3669; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3671 = 8'h44 == _io_out_bits_T_13 ? arr_68 : _GEN_3670; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3672 = 8'h45 == _io_out_bits_T_13 ? arr_69 : _GEN_3671; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3673 = 8'h46 == _io_out_bits_T_13 ? arr_70 : _GEN_3672; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3674 = 8'h47 == _io_out_bits_T_13 ? arr_71 : _GEN_3673; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3675 = 8'h48 == _io_out_bits_T_13 ? arr_72 : _GEN_3674; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3676 = 8'h49 == _io_out_bits_T_13 ? arr_73 : _GEN_3675; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3677 = 8'h4a == _io_out_bits_T_13 ? arr_74 : _GEN_3676; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3678 = 8'h4b == _io_out_bits_T_13 ? arr_75 : _GEN_3677; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3679 = 8'h4c == _io_out_bits_T_13 ? arr_76 : _GEN_3678; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3680 = 8'h4d == _io_out_bits_T_13 ? arr_77 : _GEN_3679; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3681 = 8'h4e == _io_out_bits_T_13 ? arr_78 : _GEN_3680; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3682 = 8'h4f == _io_out_bits_T_13 ? arr_79 : _GEN_3681; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3683 = 8'h50 == _io_out_bits_T_13 ? arr_80 : _GEN_3682; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3684 = 8'h51 == _io_out_bits_T_13 ? arr_81 : _GEN_3683; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3685 = 8'h52 == _io_out_bits_T_13 ? arr_82 : _GEN_3684; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3686 = 8'h53 == _io_out_bits_T_13 ? arr_83 : _GEN_3685; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3687 = 8'h54 == _io_out_bits_T_13 ? arr_84 : _GEN_3686; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3688 = 8'h55 == _io_out_bits_T_13 ? arr_85 : _GEN_3687; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3689 = 8'h56 == _io_out_bits_T_13 ? arr_86 : _GEN_3688; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3690 = 8'h57 == _io_out_bits_T_13 ? arr_87 : _GEN_3689; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3691 = 8'h58 == _io_out_bits_T_13 ? arr_88 : _GEN_3690; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3692 = 8'h59 == _io_out_bits_T_13 ? arr_89 : _GEN_3691; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3693 = 8'h5a == _io_out_bits_T_13 ? arr_90 : _GEN_3692; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3694 = 8'h5b == _io_out_bits_T_13 ? arr_91 : _GEN_3693; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3695 = 8'h5c == _io_out_bits_T_13 ? arr_92 : _GEN_3694; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3696 = 8'h5d == _io_out_bits_T_13 ? arr_93 : _GEN_3695; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3697 = 8'h5e == _io_out_bits_T_13 ? arr_94 : _GEN_3696; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3698 = 8'h5f == _io_out_bits_T_13 ? arr_95 : _GEN_3697; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3699 = 8'h60 == _io_out_bits_T_13 ? arr_96 : _GEN_3698; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3700 = 8'h61 == _io_out_bits_T_13 ? arr_97 : _GEN_3699; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3701 = 8'h62 == _io_out_bits_T_13 ? arr_98 : _GEN_3700; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3702 = 8'h63 == _io_out_bits_T_13 ? arr_99 : _GEN_3701; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3703 = 8'h64 == _io_out_bits_T_13 ? arr_100 : _GEN_3702; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3704 = 8'h65 == _io_out_bits_T_13 ? arr_101 : _GEN_3703; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3705 = 8'h66 == _io_out_bits_T_13 ? arr_102 : _GEN_3704; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3706 = 8'h67 == _io_out_bits_T_13 ? arr_103 : _GEN_3705; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3707 = 8'h68 == _io_out_bits_T_13 ? arr_104 : _GEN_3706; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3708 = 8'h69 == _io_out_bits_T_13 ? arr_105 : _GEN_3707; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3709 = 8'h6a == _io_out_bits_T_13 ? arr_106 : _GEN_3708; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3710 = 8'h6b == _io_out_bits_T_13 ? arr_107 : _GEN_3709; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3711 = 8'h6c == _io_out_bits_T_13 ? arr_108 : _GEN_3710; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3712 = 8'h6d == _io_out_bits_T_13 ? arr_109 : _GEN_3711; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3713 = 8'h6e == _io_out_bits_T_13 ? arr_110 : _GEN_3712; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3714 = 8'h6f == _io_out_bits_T_13 ? arr_111 : _GEN_3713; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3715 = 8'h70 == _io_out_bits_T_13 ? arr_112 : _GEN_3714; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3716 = 8'h71 == _io_out_bits_T_13 ? arr_113 : _GEN_3715; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3717 = 8'h72 == _io_out_bits_T_13 ? arr_114 : _GEN_3716; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3718 = 8'h73 == _io_out_bits_T_13 ? arr_115 : _GEN_3717; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3719 = 8'h74 == _io_out_bits_T_13 ? arr_116 : _GEN_3718; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3720 = 8'h75 == _io_out_bits_T_13 ? arr_117 : _GEN_3719; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3721 = 8'h76 == _io_out_bits_T_13 ? arr_118 : _GEN_3720; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3722 = 8'h77 == _io_out_bits_T_13 ? arr_119 : _GEN_3721; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3723 = 8'h78 == _io_out_bits_T_13 ? arr_120 : _GEN_3722; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3724 = 8'h79 == _io_out_bits_T_13 ? arr_121 : _GEN_3723; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3725 = 8'h7a == _io_out_bits_T_13 ? arr_122 : _GEN_3724; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3726 = 8'h7b == _io_out_bits_T_13 ? arr_123 : _GEN_3725; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3727 = 8'h7c == _io_out_bits_T_13 ? arr_124 : _GEN_3726; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3728 = 8'h7d == _io_out_bits_T_13 ? arr_125 : _GEN_3727; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3729 = 8'h7e == _io_out_bits_T_13 ? arr_126 : _GEN_3728; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3730 = 8'h7f == _io_out_bits_T_13 ? arr_127 : _GEN_3729; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3731 = 8'h80 == _io_out_bits_T_13 ? arr_128 : _GEN_3730; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3732 = 8'h81 == _io_out_bits_T_13 ? arr_129 : _GEN_3731; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3733 = 8'h82 == _io_out_bits_T_13 ? arr_130 : _GEN_3732; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3734 = 8'h83 == _io_out_bits_T_13 ? arr_131 : _GEN_3733; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3735 = 8'h84 == _io_out_bits_T_13 ? arr_132 : _GEN_3734; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3736 = 8'h85 == _io_out_bits_T_13 ? arr_133 : _GEN_3735; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3737 = 8'h86 == _io_out_bits_T_13 ? arr_134 : _GEN_3736; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3738 = 8'h87 == _io_out_bits_T_13 ? arr_135 : _GEN_3737; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3739 = 8'h88 == _io_out_bits_T_13 ? arr_136 : _GEN_3738; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3740 = 8'h89 == _io_out_bits_T_13 ? arr_137 : _GEN_3739; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3741 = 8'h8a == _io_out_bits_T_13 ? arr_138 : _GEN_3740; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3742 = 8'h8b == _io_out_bits_T_13 ? arr_139 : _GEN_3741; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3743 = 8'h8c == _io_out_bits_T_13 ? arr_140 : _GEN_3742; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3744 = 8'h8d == _io_out_bits_T_13 ? arr_141 : _GEN_3743; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3745 = 8'h8e == _io_out_bits_T_13 ? arr_142 : _GEN_3744; // @[Cat.scala 31:{58,58}]
  wire [7:0] _GEN_3746 = 8'h8f == _io_out_bits_T_13 ? arr_143 : _GEN_3745; // @[Cat.scala 31:{58,58}]
  wire [39:0] io_out_bits_hi = {_GEN_3458,_GEN_3602,_GEN_3746,_GEN_3170,_GEN_3314}; // @[Cat.scala 31:58]
  assign io_in_ready = ~full; // @[WidthConverter.scala 79:20]
  assign io_out_valid = ~empty; // @[WidthConverter.scala 80:21]
  assign io_out_bits = {io_out_bits_hi,io_out_bits_lo}; // @[Cat.scala 31:58]
  always @(posedge clock) begin
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_0 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h0 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_0 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h0 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_0 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_0 <= _GEN_1873;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_1 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h1 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_1 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h1 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_1 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_1 <= _GEN_1874;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_2 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h2 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_2 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h2 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_2 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_2 <= _GEN_1875;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_3 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h3 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_3 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h3 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_3 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_3 <= _GEN_1876;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_4 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h4 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_4 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h4 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_4 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_4 <= _GEN_1877;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_5 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h5 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_5 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h5 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_5 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_5 <= _GEN_1878;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_6 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h6 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_6 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h6 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_6 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_6 <= _GEN_1879;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_7 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h7 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_7 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h7 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_7 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_7 <= _GEN_1880;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_8 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h8 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_8 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h8 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_8 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_8 <= _GEN_1881;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_9 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h9 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_9 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h9 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_9 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_9 <= _GEN_1882;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_10 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'ha == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_10 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'ha == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_10 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_10 <= _GEN_1883;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_11 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'hb == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_11 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'hb == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_11 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_11 <= _GEN_1884;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_12 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'hc == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_12 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'hc == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_12 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_12 <= _GEN_1885;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_13 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'hd == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_13 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'hd == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_13 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_13 <= _GEN_1886;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_14 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'he == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_14 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'he == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_14 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_14 <= _GEN_1887;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_15 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'hf == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_15 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'hf == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_15 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_15 <= _GEN_1888;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_16 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h10 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_16 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h10 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_16 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_16 <= _GEN_1889;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_17 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h11 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_17 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h11 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_17 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_17 <= _GEN_1890;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_18 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h12 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_18 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h12 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_18 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_18 <= _GEN_1891;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_19 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h13 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_19 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h13 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_19 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_19 <= _GEN_1892;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_20 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h14 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_20 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h14 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_20 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_20 <= _GEN_1893;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_21 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h15 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_21 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h15 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_21 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_21 <= _GEN_1894;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_22 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h16 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_22 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h16 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_22 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_22 <= _GEN_1895;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_23 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h17 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_23 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h17 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_23 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_23 <= _GEN_1896;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_24 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h18 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_24 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h18 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_24 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_24 <= _GEN_1897;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_25 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h19 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_25 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h19 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_25 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_25 <= _GEN_1898;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_26 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h1a == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_26 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h1a == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_26 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_26 <= _GEN_1899;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_27 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h1b == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_27 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h1b == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_27 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_27 <= _GEN_1900;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_28 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h1c == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_28 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h1c == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_28 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_28 <= _GEN_1901;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_29 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h1d == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_29 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h1d == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_29 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_29 <= _GEN_1902;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_30 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h1e == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_30 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h1e == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_30 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_30 <= _GEN_1903;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_31 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h1f == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_31 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h1f == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_31 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_31 <= _GEN_1904;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_32 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h20 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_32 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h20 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_32 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_32 <= _GEN_1905;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_33 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h21 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_33 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h21 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_33 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_33 <= _GEN_1906;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_34 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h22 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_34 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h22 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_34 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_34 <= _GEN_1907;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_35 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h23 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_35 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h23 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_35 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_35 <= _GEN_1908;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_36 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h24 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_36 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h24 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_36 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_36 <= _GEN_1909;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_37 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h25 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_37 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h25 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_37 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_37 <= _GEN_1910;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_38 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h26 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_38 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h26 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_38 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_38 <= _GEN_1911;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_39 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h27 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_39 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h27 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_39 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_39 <= _GEN_1912;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_40 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h28 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_40 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h28 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_40 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_40 <= _GEN_1913;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_41 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h29 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_41 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h29 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_41 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_41 <= _GEN_1914;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_42 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h2a == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_42 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h2a == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_42 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_42 <= _GEN_1915;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_43 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h2b == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_43 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h2b == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_43 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_43 <= _GEN_1916;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_44 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h2c == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_44 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h2c == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_44 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_44 <= _GEN_1917;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_45 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h2d == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_45 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h2d == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_45 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_45 <= _GEN_1918;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_46 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h2e == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_46 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h2e == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_46 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_46 <= _GEN_1919;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_47 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h2f == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_47 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h2f == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_47 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_47 <= _GEN_1920;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_48 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h30 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_48 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h30 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_48 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_48 <= _GEN_1921;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_49 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h31 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_49 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h31 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_49 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_49 <= _GEN_1922;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_50 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h32 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_50 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h32 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_50 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_50 <= _GEN_1923;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_51 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h33 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_51 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h33 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_51 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_51 <= _GEN_1924;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_52 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h34 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_52 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h34 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_52 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_52 <= _GEN_1925;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_53 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h35 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_53 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h35 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_53 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_53 <= _GEN_1926;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_54 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h36 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_54 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h36 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_54 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_54 <= _GEN_1927;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_55 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h37 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_55 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h37 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_55 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_55 <= _GEN_1928;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_56 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h38 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_56 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h38 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_56 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_56 <= _GEN_1929;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_57 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h39 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_57 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h39 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_57 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_57 <= _GEN_1930;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_58 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h3a == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_58 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h3a == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_58 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_58 <= _GEN_1931;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_59 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h3b == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_59 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h3b == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_59 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_59 <= _GEN_1932;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_60 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h3c == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_60 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h3c == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_60 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_60 <= _GEN_1933;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_61 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h3d == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_61 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h3d == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_61 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_61 <= _GEN_1934;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_62 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h3e == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_62 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h3e == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_62 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_62 <= _GEN_1935;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_63 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h3f == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_63 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h3f == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_63 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_63 <= _GEN_1936;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_64 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h40 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_64 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h40 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_64 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_64 <= _GEN_1937;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_65 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h41 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_65 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h41 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_65 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_65 <= _GEN_1938;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_66 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h42 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_66 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h42 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_66 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_66 <= _GEN_1939;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_67 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h43 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_67 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h43 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_67 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_67 <= _GEN_1940;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_68 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h44 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_68 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h44 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_68 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_68 <= _GEN_1941;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_69 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h45 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_69 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h45 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_69 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_69 <= _GEN_1942;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_70 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h46 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_70 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h46 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_70 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_70 <= _GEN_1943;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_71 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h47 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_71 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h47 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_71 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_71 <= _GEN_1944;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_72 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h48 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_72 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h48 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_72 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_72 <= _GEN_1945;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_73 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h49 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_73 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h49 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_73 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_73 <= _GEN_1946;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_74 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h4a == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_74 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h4a == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_74 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_74 <= _GEN_1947;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_75 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h4b == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_75 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h4b == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_75 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_75 <= _GEN_1948;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_76 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h4c == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_76 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h4c == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_76 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_76 <= _GEN_1949;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_77 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h4d == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_77 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h4d == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_77 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_77 <= _GEN_1950;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_78 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h4e == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_78 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h4e == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_78 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_78 <= _GEN_1951;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_79 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h4f == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_79 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h4f == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_79 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_79 <= _GEN_1952;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_80 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h50 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_80 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h50 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_80 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_80 <= _GEN_1953;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_81 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h51 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_81 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h51 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_81 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_81 <= _GEN_1954;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_82 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h52 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_82 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h52 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_82 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_82 <= _GEN_1955;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_83 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h53 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_83 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h53 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_83 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_83 <= _GEN_1956;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_84 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h54 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_84 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h54 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_84 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_84 <= _GEN_1957;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_85 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h55 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_85 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h55 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_85 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_85 <= _GEN_1958;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_86 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h56 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_86 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h56 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_86 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_86 <= _GEN_1959;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_87 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h57 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_87 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h57 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_87 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_87 <= _GEN_1960;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_88 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h58 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_88 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h58 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_88 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_88 <= _GEN_1961;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_89 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h59 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_89 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h59 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_89 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_89 <= _GEN_1962;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_90 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h5a == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_90 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h5a == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_90 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_90 <= _GEN_1963;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_91 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h5b == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_91 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h5b == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_91 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_91 <= _GEN_1964;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_92 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h5c == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_92 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h5c == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_92 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_92 <= _GEN_1965;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_93 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h5d == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_93 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h5d == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_93 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_93 <= _GEN_1966;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_94 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h5e == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_94 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h5e == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_94 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_94 <= _GEN_1967;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_95 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h5f == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_95 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h5f == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_95 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_95 <= _GEN_1968;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_96 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h60 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_96 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h60 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_96 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_96 <= _GEN_1969;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_97 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h61 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_97 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h61 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_97 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_97 <= _GEN_1970;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_98 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h62 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_98 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h62 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_98 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_98 <= _GEN_1971;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_99 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h63 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_99 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h63 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_99 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_99 <= _GEN_1972;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_100 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h64 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_100 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h64 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_100 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_100 <= _GEN_1973;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_101 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h65 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_101 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h65 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_101 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_101 <= _GEN_1974;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_102 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h66 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_102 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h66 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_102 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_102 <= _GEN_1975;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_103 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h67 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_103 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h67 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_103 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_103 <= _GEN_1976;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_104 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h68 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_104 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h68 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_104 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_104 <= _GEN_1977;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_105 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h69 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_105 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h69 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_105 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_105 <= _GEN_1978;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_106 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h6a == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_106 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h6a == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_106 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_106 <= _GEN_1979;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_107 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h6b == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_107 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h6b == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_107 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_107 <= _GEN_1980;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_108 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h6c == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_108 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h6c == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_108 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_108 <= _GEN_1981;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_109 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h6d == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_109 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h6d == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_109 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_109 <= _GEN_1982;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_110 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h6e == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_110 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h6e == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_110 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_110 <= _GEN_1983;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_111 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h6f == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_111 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h6f == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_111 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_111 <= _GEN_1984;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_112 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h70 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_112 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h70 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_112 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_112 <= _GEN_1985;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_113 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h71 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_113 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h71 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_113 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_113 <= _GEN_1986;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_114 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h72 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_114 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h72 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_114 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_114 <= _GEN_1987;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_115 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h73 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_115 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h73 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_115 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_115 <= _GEN_1988;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_116 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h74 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_116 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h74 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_116 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_116 <= _GEN_1989;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_117 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h75 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_117 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h75 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_117 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_117 <= _GEN_1990;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_118 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h76 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_118 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h76 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_118 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_118 <= _GEN_1991;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_119 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h77 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_119 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h77 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_119 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_119 <= _GEN_1992;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_120 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h78 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_120 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h78 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_120 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_120 <= _GEN_1993;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_121 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h79 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_121 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h79 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_121 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_121 <= _GEN_1994;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_122 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h7a == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_122 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h7a == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_122 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_122 <= _GEN_1995;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_123 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h7b == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_123 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h7b == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_123 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_123 <= _GEN_1996;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_124 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h7c == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_124 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h7c == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_124 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_124 <= _GEN_1997;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_125 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h7d == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_125 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h7d == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_125 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_125 <= _GEN_1998;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_126 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h7e == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_126 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h7e == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_126 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_126 <= _GEN_1999;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_127 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h7f == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_127 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h7f == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_127 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_127 <= _GEN_2000;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_128 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h80 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_128 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h80 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_128 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_128 <= _GEN_2001;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_129 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h81 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_129 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h81 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_129 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_129 <= _GEN_2002;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_130 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h82 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_130 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h82 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_130 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_130 <= _GEN_2003;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_131 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h83 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_131 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h83 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_131 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_131 <= _GEN_2004;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_132 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h84 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_132 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h84 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_132 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_132 <= _GEN_2005;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_133 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h85 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_133 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h85 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_133 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_133 <= _GEN_2006;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_134 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h86 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_134 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h86 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_134 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_134 <= _GEN_2007;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_135 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h87 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_135 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h87 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_135 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_135 <= _GEN_2008;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_136 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h88 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_136 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h88 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_136 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_136 <= _GEN_2009;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_137 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h89 == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_137 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h89 == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_137 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_137 <= _GEN_2010;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_138 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h8a == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_138 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h8a == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_138 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_138 <= _GEN_2011;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_139 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h8b == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_139 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h8b == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_139 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_139 <= _GEN_2012;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_140 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h8c == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_140 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h8c == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_140 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_140 <= _GEN_2013;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_141 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h8d == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_141 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h8d == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_141 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_141 <= _GEN_2014;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_142 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h8e == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_142 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h8e == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_142 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_142 <= _GEN_2015;
      end
    end
    if (reset) begin // @[WidthConverter.scala 24:29]
      arr_143 <= 8'h0; // @[WidthConverter.scala 24:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      if (8'h8f == _T_32) begin // @[WidthConverter.scala 67:27]
        arr_143 <= io_in_bits[127:120]; // @[WidthConverter.scala 67:27]
      end else if (8'h8f == _T_30) begin // @[WidthConverter.scala 67:27]
        arr_143 <= io_in_bits[119:112]; // @[WidthConverter.scala 67:27]
      end else begin
        arr_143 <= _GEN_2016;
      end
    end
    if (reset) begin // @[WidthConverter.scala 25:29]
      enqPtr <= 8'h0; // @[WidthConverter.scala 25:29]
    end else if (doEnq) begin // @[WidthConverter.scala 65:17]
      enqPtr <= _enqPtr_T_2; // @[WidthConverter.scala 89:9]
    end
    if (reset) begin // @[WidthConverter.scala 26:29]
      deqPtr <= 8'h0; // @[WidthConverter.scala 26:29]
    end else if (doDeq) begin // @[WidthConverter.scala 75:17]
      deqPtr <= _deqPtr_T_2; // @[WidthConverter.scala 89:9]
    end
    if (reset) begin // @[WidthConverter.scala 27:29]
      maybeFull <= 1'h0; // @[WidthConverter.scala 27:29]
    end else if (doEnq != doDeq) begin // @[WidthConverter.scala 61:27]
      maybeFull <= doEnq; // @[WidthConverter.scala 62:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  arr_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  arr_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  arr_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  arr_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  arr_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  arr_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  arr_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  arr_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  arr_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  arr_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  arr_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  arr_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  arr_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  arr_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  arr_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  arr_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  arr_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  arr_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  arr_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  arr_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  arr_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  arr_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  arr_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  arr_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  arr_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  arr_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  arr_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  arr_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  arr_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  arr_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  arr_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  arr_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  arr_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  arr_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  arr_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  arr_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  arr_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  arr_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  arr_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  arr_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  arr_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  arr_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  arr_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  arr_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  arr_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  arr_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  arr_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  arr_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  arr_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  arr_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  arr_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  arr_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  arr_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  arr_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  arr_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  arr_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  arr_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  arr_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  arr_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  arr_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  arr_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  arr_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  arr_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  arr_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  arr_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  arr_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  arr_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  arr_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  arr_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  arr_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  arr_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  arr_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  arr_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  arr_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  arr_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  arr_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  arr_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  arr_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  arr_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  arr_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  arr_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  arr_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  arr_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  arr_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  arr_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  arr_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  arr_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  arr_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  arr_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  arr_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  arr_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  arr_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  arr_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  arr_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  arr_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  arr_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  arr_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  arr_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  arr_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  arr_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  arr_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  arr_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  arr_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  arr_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  arr_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  arr_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  arr_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  arr_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  arr_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  arr_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  arr_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  arr_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  arr_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  arr_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  arr_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  arr_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  arr_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  arr_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  arr_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  arr_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  arr_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  arr_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  arr_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  arr_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  arr_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  arr_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  arr_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  arr_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  arr_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  arr_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  arr_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  arr_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  arr_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  arr_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  arr_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  arr_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  arr_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  arr_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  arr_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  arr_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  arr_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  arr_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  arr_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  arr_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  enqPtr = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  deqPtr = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  maybeFull = _RAND_146[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Transmission(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits,
  input          io_out_ready,
  output         io_out_valid,
  output [71:0]  io_out_bits
);
  wire  widthConverter_clock; // @[Transmission.scala 19:32]
  wire  widthConverter_reset; // @[Transmission.scala 19:32]
  wire  widthConverter_io_in_ready; // @[Transmission.scala 19:32]
  wire  widthConverter_io_in_valid; // @[Transmission.scala 19:32]
  wire [127:0] widthConverter_io_in_bits; // @[Transmission.scala 19:32]
  wire  widthConverter_io_out_ready; // @[Transmission.scala 19:32]
  wire  widthConverter_io_out_valid; // @[Transmission.scala 19:32]
  wire [71:0] widthConverter_io_out_bits; // @[Transmission.scala 19:32]
  WidthConverter widthConverter ( // @[Transmission.scala 19:32]
    .clock(widthConverter_clock),
    .reset(widthConverter_reset),
    .io_in_ready(widthConverter_io_in_ready),
    .io_in_valid(widthConverter_io_in_valid),
    .io_in_bits(widthConverter_io_in_bits),
    .io_out_ready(widthConverter_io_out_ready),
    .io_out_valid(widthConverter_io_out_valid),
    .io_out_bits(widthConverter_io_out_bits)
  );
  assign io_in_ready = widthConverter_io_in_ready; // @[Transmission.scala 20:26]
  assign io_out_valid = widthConverter_io_out_valid; // @[Transmission.scala 21:12]
  assign io_out_bits = widthConverter_io_out_bits; // @[Transmission.scala 21:12]
  assign widthConverter_clock = clock;
  assign widthConverter_reset = reset;
  assign widthConverter_io_in_valid = io_in_valid; // @[Transmission.scala 20:26]
  assign widthConverter_io_in_bits = io_in_bits; // @[Transmission.scala 20:26]
  assign widthConverter_io_out_ready = io_out_ready; // @[Transmission.scala 21:12]
endmodule
module top_zcu104(
  input          clock,
  input          reset,
  input  [127:0] instruction_tdata,
  input          instruction_tvalid,
  output         instruction_tready,
  input          instruction_tlast,
  input          m_axi_dram0_awready,
  output         m_axi_dram0_awvalid,
  output [5:0]   m_axi_dram0_awid,
  output [31:0]  m_axi_dram0_awaddr,
  output [7:0]   m_axi_dram0_awlen,
  output [2:0]   m_axi_dram0_awsize,
  output [1:0]   m_axi_dram0_awburst,
  output [1:0]   m_axi_dram0_awlock,
  output [3:0]   m_axi_dram0_awcache,
  output [2:0]   m_axi_dram0_awprot,
  output [3:0]   m_axi_dram0_awqos,
  input          m_axi_dram0_wready,
  output         m_axi_dram0_wvalid,
  output [5:0]   m_axi_dram0_wid,
  output [127:0] m_axi_dram0_wdata,
  output [15:0]  m_axi_dram0_wstrb,
  output         m_axi_dram0_wlast,
  output         m_axi_dram0_bready,
  input          m_axi_dram0_bvalid,
  input  [5:0]   m_axi_dram0_bid,
  input  [1:0]   m_axi_dram0_bresp,
  input          m_axi_dram0_arready,
  output         m_axi_dram0_arvalid,
  output [5:0]   m_axi_dram0_arid,
  output [31:0]  m_axi_dram0_araddr,
  output [7:0]   m_axi_dram0_arlen,
  output [2:0]   m_axi_dram0_arsize,
  output [1:0]   m_axi_dram0_arburst,
  output [1:0]   m_axi_dram0_arlock,
  output [3:0]   m_axi_dram0_arcache,
  output [2:0]   m_axi_dram0_arprot,
  output [3:0]   m_axi_dram0_arqos,
  output         m_axi_dram0_rready,
  input          m_axi_dram0_rvalid,
  input  [5:0]   m_axi_dram0_rid,
  input  [127:0] m_axi_dram0_rdata,
  input  [1:0]   m_axi_dram0_rresp,
  input          m_axi_dram0_rlast,
  input          m_axi_dram1_awready,
  output         m_axi_dram1_awvalid,
  output [5:0]   m_axi_dram1_awid,
  output [31:0]  m_axi_dram1_awaddr,
  output [7:0]   m_axi_dram1_awlen,
  output [2:0]   m_axi_dram1_awsize,
  output [1:0]   m_axi_dram1_awburst,
  output [1:0]   m_axi_dram1_awlock,
  output [3:0]   m_axi_dram1_awcache,
  output [2:0]   m_axi_dram1_awprot,
  output [3:0]   m_axi_dram1_awqos,
  input          m_axi_dram1_wready,
  output         m_axi_dram1_wvalid,
  output [5:0]   m_axi_dram1_wid,
  output [127:0] m_axi_dram1_wdata,
  output [15:0]  m_axi_dram1_wstrb,
  output         m_axi_dram1_wlast,
  output         m_axi_dram1_bready,
  input          m_axi_dram1_bvalid,
  input  [5:0]   m_axi_dram1_bid,
  input  [1:0]   m_axi_dram1_bresp,
  input          m_axi_dram1_arready,
  output         m_axi_dram1_arvalid,
  output [5:0]   m_axi_dram1_arid,
  output [31:0]  m_axi_dram1_araddr,
  output [7:0]   m_axi_dram1_arlen,
  output [2:0]   m_axi_dram1_arsize,
  output [1:0]   m_axi_dram1_arburst,
  output [1:0]   m_axi_dram1_arlock,
  output [3:0]   m_axi_dram1_arcache,
  output [2:0]   m_axi_dram1_arprot,
  output [3:0]   m_axi_dram1_arqos,
  output         m_axi_dram1_rready,
  input          m_axi_dram1_rvalid,
  input  [5:0]   m_axi_dram1_rid,
  input  [127:0] m_axi_dram1_rdata,
  input  [1:0]   m_axi_dram1_rresp,
  input          m_axi_dram1_rlast
);
  wire  tcu_clock; // @[Top.scala 76:21]
  wire  tcu_reset; // @[Top.scala 76:21]
  wire  tcu_instruction_ready; // @[Top.scala 76:21]
  wire  tcu_instruction_valid; // @[Top.scala 76:21]
  wire [3:0] tcu_instruction_bits_opcode; // @[Top.scala 76:21]
  wire [3:0] tcu_instruction_bits_flags; // @[Top.scala 76:21]
  wire [63:0] tcu_instruction_bits_arguments; // @[Top.scala 76:21]
  wire  tcu_dram0_writeAddress_ready; // @[Top.scala 76:21]
  wire  tcu_dram0_writeAddress_valid; // @[Top.scala 76:21]
  wire [5:0] tcu_dram0_writeAddress_bits_id; // @[Top.scala 76:21]
  wire [31:0] tcu_dram0_writeAddress_bits_addr; // @[Top.scala 76:21]
  wire [7:0] tcu_dram0_writeAddress_bits_len; // @[Top.scala 76:21]
  wire [2:0] tcu_dram0_writeAddress_bits_size; // @[Top.scala 76:21]
  wire [1:0] tcu_dram0_writeAddress_bits_burst; // @[Top.scala 76:21]
  wire [1:0] tcu_dram0_writeAddress_bits_lock; // @[Top.scala 76:21]
  wire [3:0] tcu_dram0_writeAddress_bits_cache; // @[Top.scala 76:21]
  wire [2:0] tcu_dram0_writeAddress_bits_prot; // @[Top.scala 76:21]
  wire [3:0] tcu_dram0_writeAddress_bits_qos; // @[Top.scala 76:21]
  wire  tcu_dram0_writeData_ready; // @[Top.scala 76:21]
  wire  tcu_dram0_writeData_valid; // @[Top.scala 76:21]
  wire [5:0] tcu_dram0_writeData_bits_id; // @[Top.scala 76:21]
  wire [127:0] tcu_dram0_writeData_bits_data; // @[Top.scala 76:21]
  wire [15:0] tcu_dram0_writeData_bits_strb; // @[Top.scala 76:21]
  wire  tcu_dram0_writeData_bits_last; // @[Top.scala 76:21]
  wire  tcu_dram0_writeResponse_ready; // @[Top.scala 76:21]
  wire  tcu_dram0_writeResponse_valid; // @[Top.scala 76:21]
  wire  tcu_dram0_readAddress_ready; // @[Top.scala 76:21]
  wire  tcu_dram0_readAddress_valid; // @[Top.scala 76:21]
  wire [5:0] tcu_dram0_readAddress_bits_id; // @[Top.scala 76:21]
  wire [31:0] tcu_dram0_readAddress_bits_addr; // @[Top.scala 76:21]
  wire [7:0] tcu_dram0_readAddress_bits_len; // @[Top.scala 76:21]
  wire [2:0] tcu_dram0_readAddress_bits_size; // @[Top.scala 76:21]
  wire [1:0] tcu_dram0_readAddress_bits_burst; // @[Top.scala 76:21]
  wire [1:0] tcu_dram0_readAddress_bits_lock; // @[Top.scala 76:21]
  wire [3:0] tcu_dram0_readAddress_bits_cache; // @[Top.scala 76:21]
  wire [2:0] tcu_dram0_readAddress_bits_prot; // @[Top.scala 76:21]
  wire [3:0] tcu_dram0_readAddress_bits_qos; // @[Top.scala 76:21]
  wire  tcu_dram0_readData_ready; // @[Top.scala 76:21]
  wire  tcu_dram0_readData_valid; // @[Top.scala 76:21]
  wire [127:0] tcu_dram0_readData_bits_data; // @[Top.scala 76:21]
  wire  tcu_dram1_writeAddress_ready; // @[Top.scala 76:21]
  wire  tcu_dram1_writeAddress_valid; // @[Top.scala 76:21]
  wire [5:0] tcu_dram1_writeAddress_bits_id; // @[Top.scala 76:21]
  wire [31:0] tcu_dram1_writeAddress_bits_addr; // @[Top.scala 76:21]
  wire [7:0] tcu_dram1_writeAddress_bits_len; // @[Top.scala 76:21]
  wire [2:0] tcu_dram1_writeAddress_bits_size; // @[Top.scala 76:21]
  wire [1:0] tcu_dram1_writeAddress_bits_burst; // @[Top.scala 76:21]
  wire [1:0] tcu_dram1_writeAddress_bits_lock; // @[Top.scala 76:21]
  wire [3:0] tcu_dram1_writeAddress_bits_cache; // @[Top.scala 76:21]
  wire [2:0] tcu_dram1_writeAddress_bits_prot; // @[Top.scala 76:21]
  wire [3:0] tcu_dram1_writeAddress_bits_qos; // @[Top.scala 76:21]
  wire  tcu_dram1_writeData_ready; // @[Top.scala 76:21]
  wire  tcu_dram1_writeData_valid; // @[Top.scala 76:21]
  wire [5:0] tcu_dram1_writeData_bits_id; // @[Top.scala 76:21]
  wire [127:0] tcu_dram1_writeData_bits_data; // @[Top.scala 76:21]
  wire [15:0] tcu_dram1_writeData_bits_strb; // @[Top.scala 76:21]
  wire  tcu_dram1_writeData_bits_last; // @[Top.scala 76:21]
  wire  tcu_dram1_writeResponse_ready; // @[Top.scala 76:21]
  wire  tcu_dram1_writeResponse_valid; // @[Top.scala 76:21]
  wire  tcu_dram1_readAddress_ready; // @[Top.scala 76:21]
  wire  tcu_dram1_readAddress_valid; // @[Top.scala 76:21]
  wire [5:0] tcu_dram1_readAddress_bits_id; // @[Top.scala 76:21]
  wire [31:0] tcu_dram1_readAddress_bits_addr; // @[Top.scala 76:21]
  wire [7:0] tcu_dram1_readAddress_bits_len; // @[Top.scala 76:21]
  wire [2:0] tcu_dram1_readAddress_bits_size; // @[Top.scala 76:21]
  wire [1:0] tcu_dram1_readAddress_bits_burst; // @[Top.scala 76:21]
  wire [1:0] tcu_dram1_readAddress_bits_lock; // @[Top.scala 76:21]
  wire [3:0] tcu_dram1_readAddress_bits_cache; // @[Top.scala 76:21]
  wire [2:0] tcu_dram1_readAddress_bits_prot; // @[Top.scala 76:21]
  wire [3:0] tcu_dram1_readAddress_bits_qos; // @[Top.scala 76:21]
  wire  tcu_dram1_readData_ready; // @[Top.scala 76:21]
  wire  tcu_dram1_readData_valid; // @[Top.scala 76:21]
  wire [127:0] tcu_dram1_readData_bits_data; // @[Top.scala 76:21]
  wire  transmission_clock; // @[package.scala 27:30]
  wire  transmission_reset; // @[package.scala 27:30]
  wire  transmission_io_in_ready; // @[package.scala 27:30]
  wire  transmission_io_in_valid; // @[package.scala 27:30]
  wire [127:0] transmission_io_in_bits; // @[package.scala 27:30]
  wire  transmission_io_out_ready; // @[package.scala 27:30]
  wire  transmission_io_out_valid; // @[package.scala 27:30]
  wire [71:0] transmission_io_out_bits; // @[package.scala 27:30]
  wire [71:0] _tcu_instruction_bits_WIRE_1 = transmission_io_out_bits;
  AXIWrapperTCU tcu ( // @[Top.scala 76:21]
    .clock(tcu_clock),
    .reset(tcu_reset),
    .instruction_ready(tcu_instruction_ready),
    .instruction_valid(tcu_instruction_valid),
    .instruction_bits_opcode(tcu_instruction_bits_opcode),
    .instruction_bits_flags(tcu_instruction_bits_flags),
    .instruction_bits_arguments(tcu_instruction_bits_arguments),
    .dram0_writeAddress_ready(tcu_dram0_writeAddress_ready),
    .dram0_writeAddress_valid(tcu_dram0_writeAddress_valid),
    .dram0_writeAddress_bits_id(tcu_dram0_writeAddress_bits_id),
    .dram0_writeAddress_bits_addr(tcu_dram0_writeAddress_bits_addr),
    .dram0_writeAddress_bits_len(tcu_dram0_writeAddress_bits_len),
    .dram0_writeAddress_bits_size(tcu_dram0_writeAddress_bits_size),
    .dram0_writeAddress_bits_burst(tcu_dram0_writeAddress_bits_burst),
    .dram0_writeAddress_bits_lock(tcu_dram0_writeAddress_bits_lock),
    .dram0_writeAddress_bits_cache(tcu_dram0_writeAddress_bits_cache),
    .dram0_writeAddress_bits_prot(tcu_dram0_writeAddress_bits_prot),
    .dram0_writeAddress_bits_qos(tcu_dram0_writeAddress_bits_qos),
    .dram0_writeData_ready(tcu_dram0_writeData_ready),
    .dram0_writeData_valid(tcu_dram0_writeData_valid),
    .dram0_writeData_bits_id(tcu_dram0_writeData_bits_id),
    .dram0_writeData_bits_data(tcu_dram0_writeData_bits_data),
    .dram0_writeData_bits_strb(tcu_dram0_writeData_bits_strb),
    .dram0_writeData_bits_last(tcu_dram0_writeData_bits_last),
    .dram0_writeResponse_ready(tcu_dram0_writeResponse_ready),
    .dram0_writeResponse_valid(tcu_dram0_writeResponse_valid),
    .dram0_readAddress_ready(tcu_dram0_readAddress_ready),
    .dram0_readAddress_valid(tcu_dram0_readAddress_valid),
    .dram0_readAddress_bits_id(tcu_dram0_readAddress_bits_id),
    .dram0_readAddress_bits_addr(tcu_dram0_readAddress_bits_addr),
    .dram0_readAddress_bits_len(tcu_dram0_readAddress_bits_len),
    .dram0_readAddress_bits_size(tcu_dram0_readAddress_bits_size),
    .dram0_readAddress_bits_burst(tcu_dram0_readAddress_bits_burst),
    .dram0_readAddress_bits_lock(tcu_dram0_readAddress_bits_lock),
    .dram0_readAddress_bits_cache(tcu_dram0_readAddress_bits_cache),
    .dram0_readAddress_bits_prot(tcu_dram0_readAddress_bits_prot),
    .dram0_readAddress_bits_qos(tcu_dram0_readAddress_bits_qos),
    .dram0_readData_ready(tcu_dram0_readData_ready),
    .dram0_readData_valid(tcu_dram0_readData_valid),
    .dram0_readData_bits_data(tcu_dram0_readData_bits_data),
    .dram1_writeAddress_ready(tcu_dram1_writeAddress_ready),
    .dram1_writeAddress_valid(tcu_dram1_writeAddress_valid),
    .dram1_writeAddress_bits_id(tcu_dram1_writeAddress_bits_id),
    .dram1_writeAddress_bits_addr(tcu_dram1_writeAddress_bits_addr),
    .dram1_writeAddress_bits_len(tcu_dram1_writeAddress_bits_len),
    .dram1_writeAddress_bits_size(tcu_dram1_writeAddress_bits_size),
    .dram1_writeAddress_bits_burst(tcu_dram1_writeAddress_bits_burst),
    .dram1_writeAddress_bits_lock(tcu_dram1_writeAddress_bits_lock),
    .dram1_writeAddress_bits_cache(tcu_dram1_writeAddress_bits_cache),
    .dram1_writeAddress_bits_prot(tcu_dram1_writeAddress_bits_prot),
    .dram1_writeAddress_bits_qos(tcu_dram1_writeAddress_bits_qos),
    .dram1_writeData_ready(tcu_dram1_writeData_ready),
    .dram1_writeData_valid(tcu_dram1_writeData_valid),
    .dram1_writeData_bits_id(tcu_dram1_writeData_bits_id),
    .dram1_writeData_bits_data(tcu_dram1_writeData_bits_data),
    .dram1_writeData_bits_strb(tcu_dram1_writeData_bits_strb),
    .dram1_writeData_bits_last(tcu_dram1_writeData_bits_last),
    .dram1_writeResponse_ready(tcu_dram1_writeResponse_ready),
    .dram1_writeResponse_valid(tcu_dram1_writeResponse_valid),
    .dram1_readAddress_ready(tcu_dram1_readAddress_ready),
    .dram1_readAddress_valid(tcu_dram1_readAddress_valid),
    .dram1_readAddress_bits_id(tcu_dram1_readAddress_bits_id),
    .dram1_readAddress_bits_addr(tcu_dram1_readAddress_bits_addr),
    .dram1_readAddress_bits_len(tcu_dram1_readAddress_bits_len),
    .dram1_readAddress_bits_size(tcu_dram1_readAddress_bits_size),
    .dram1_readAddress_bits_burst(tcu_dram1_readAddress_bits_burst),
    .dram1_readAddress_bits_lock(tcu_dram1_readAddress_bits_lock),
    .dram1_readAddress_bits_cache(tcu_dram1_readAddress_bits_cache),
    .dram1_readAddress_bits_prot(tcu_dram1_readAddress_bits_prot),
    .dram1_readAddress_bits_qos(tcu_dram1_readAddress_bits_qos),
    .dram1_readData_ready(tcu_dram1_readData_ready),
    .dram1_readData_valid(tcu_dram1_readData_valid),
    .dram1_readData_bits_data(tcu_dram1_readData_bits_data)
  );
  Transmission transmission ( // @[package.scala 27:30]
    .clock(transmission_clock),
    .reset(transmission_reset),
    .io_in_ready(transmission_io_in_ready),
    .io_in_valid(transmission_io_in_valid),
    .io_in_bits(transmission_io_in_bits),
    .io_out_ready(transmission_io_out_ready),
    .io_out_valid(transmission_io_out_valid),
    .io_out_bits(transmission_io_out_bits)
  );
  assign instruction_tready = transmission_io_in_ready; // @[AXI4Stream.scala 16:17 package.scala 29:24]
  assign m_axi_dram0_awvalid = tcu_dram0_writeAddress_valid; // @[ExternalMaster.scala 68:33]
  assign m_axi_dram0_awid = tcu_dram0_writeAddress_bits_id; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_awaddr = tcu_dram0_writeAddress_bits_addr; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_awlen = tcu_dram0_writeAddress_bits_len; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_awsize = tcu_dram0_writeAddress_bits_size; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_awburst = tcu_dram0_writeAddress_bits_burst; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_awlock = tcu_dram0_writeAddress_bits_lock; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_awcache = tcu_dram0_writeAddress_bits_cache; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_awprot = tcu_dram0_writeAddress_bits_prot; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_awqos = tcu_dram0_writeAddress_bits_qos; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_wvalid = tcu_dram0_writeData_valid; // @[ExternalMaster.scala 68:33]
  assign m_axi_dram0_wid = tcu_dram0_writeData_bits_id; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_wdata = tcu_dram0_writeData_bits_data; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_wstrb = tcu_dram0_writeData_bits_strb; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_wlast = tcu_dram0_writeData_bits_last; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_bready = tcu_dram0_writeResponse_ready; // @[ExternalMaster.scala 69:33]
  assign m_axi_dram0_arvalid = tcu_dram0_readAddress_valid; // @[ExternalMaster.scala 68:33]
  assign m_axi_dram0_arid = tcu_dram0_readAddress_bits_id; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_araddr = tcu_dram0_readAddress_bits_addr; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_arlen = tcu_dram0_readAddress_bits_len; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_arsize = tcu_dram0_readAddress_bits_size; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_arburst = tcu_dram0_readAddress_bits_burst; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_arlock = tcu_dram0_readAddress_bits_lock; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_arcache = tcu_dram0_readAddress_bits_cache; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_arprot = tcu_dram0_readAddress_bits_prot; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_arqos = tcu_dram0_readAddress_bits_qos; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram0_rready = tcu_dram0_readData_ready; // @[ExternalMaster.scala 69:33]
  assign m_axi_dram1_awvalid = tcu_dram1_writeAddress_valid; // @[ExternalMaster.scala 68:33]
  assign m_axi_dram1_awid = tcu_dram1_writeAddress_bits_id; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_awaddr = tcu_dram1_writeAddress_bits_addr; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_awlen = tcu_dram1_writeAddress_bits_len; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_awsize = tcu_dram1_writeAddress_bits_size; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_awburst = tcu_dram1_writeAddress_bits_burst; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_awlock = tcu_dram1_writeAddress_bits_lock; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_awcache = tcu_dram1_writeAddress_bits_cache; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_awprot = tcu_dram1_writeAddress_bits_prot; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_awqos = tcu_dram1_writeAddress_bits_qos; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_wvalid = tcu_dram1_writeData_valid; // @[ExternalMaster.scala 68:33]
  assign m_axi_dram1_wid = tcu_dram1_writeData_bits_id; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_wdata = tcu_dram1_writeData_bits_data; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_wstrb = tcu_dram1_writeData_bits_strb; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_wlast = tcu_dram1_writeData_bits_last; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_bready = tcu_dram1_writeResponse_ready; // @[ExternalMaster.scala 69:33]
  assign m_axi_dram1_arvalid = tcu_dram1_readAddress_valid; // @[ExternalMaster.scala 68:33]
  assign m_axi_dram1_arid = tcu_dram1_readAddress_bits_id; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_araddr = tcu_dram1_readAddress_bits_addr; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_arlen = tcu_dram1_readAddress_bits_len; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_arsize = tcu_dram1_readAddress_bits_size; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_arburst = tcu_dram1_readAddress_bits_burst; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_arlock = tcu_dram1_readAddress_bits_lock; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_arcache = tcu_dram1_readAddress_bits_cache; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_arprot = tcu_dram1_readAddress_bits_prot; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_arqos = tcu_dram1_readAddress_bits_qos; // @[ExternalMaster.scala 72:26]
  assign m_axi_dram1_rready = tcu_dram1_readData_ready; // @[ExternalMaster.scala 69:33]
  assign tcu_clock = clock;
  assign tcu_reset = ~reset; // @[Top.scala 75:56]
  assign tcu_instruction_valid = transmission_io_out_valid; // @[package.scala 30:15]
  assign tcu_instruction_bits_opcode = _tcu_instruction_bits_WIRE_1[71:68]; // @[package.scala 32:50]
  assign tcu_instruction_bits_flags = _tcu_instruction_bits_WIRE_1[67:64]; // @[package.scala 32:50]
  assign tcu_instruction_bits_arguments = _tcu_instruction_bits_WIRE_1[63:0]; // @[package.scala 32:50]
  assign tcu_dram0_writeAddress_ready = m_axi_dram0_awready; // @[ExternalMaster.scala 69:33]
  assign tcu_dram0_writeData_ready = m_axi_dram0_wready; // @[ExternalMaster.scala 69:33]
  assign tcu_dram0_writeResponse_valid = m_axi_dram0_bvalid; // @[ExternalMaster.scala 68:33]
  assign tcu_dram0_readAddress_ready = m_axi_dram0_arready; // @[ExternalMaster.scala 69:33]
  assign tcu_dram0_readData_valid = m_axi_dram0_rvalid; // @[ExternalMaster.scala 68:33]
  assign tcu_dram0_readData_bits_data = m_axi_dram0_rdata; // @[ExternalMaster.scala 72:26]
  assign tcu_dram1_writeAddress_ready = m_axi_dram1_awready; // @[ExternalMaster.scala 69:33]
  assign tcu_dram1_writeData_ready = m_axi_dram1_wready; // @[ExternalMaster.scala 69:33]
  assign tcu_dram1_writeResponse_valid = m_axi_dram1_bvalid; // @[ExternalMaster.scala 68:33]
  assign tcu_dram1_readAddress_ready = m_axi_dram1_arready; // @[ExternalMaster.scala 69:33]
  assign tcu_dram1_readData_valid = m_axi_dram1_rvalid; // @[ExternalMaster.scala 68:33]
  assign tcu_dram1_readData_bits_data = m_axi_dram1_rdata; // @[ExternalMaster.scala 72:26]
  assign transmission_clock = clock;
  assign transmission_reset = ~reset; // @[Top.scala 75:56]
  assign transmission_io_in_valid = instruction_tvalid; // @[AXI4Stream.scala 16:17 18:13]
  assign transmission_io_in_bits = instruction_tdata; // @[AXI4Stream.scala 16:17 17:12]
  assign transmission_io_out_ready = tcu_instruction_ready; // @[package.scala 31:31]
endmodule
